`timescale 1ns/10ps
`include "cal1.v"
`include "cal2.v"
`define _SIZE 20
`define DECODE 0
`define ENCODE 1
`define DONE   2
module decoder # (
    parameter integer N = 1024,
    parameter integer STEP = 10,
    parameter integer SIZE = `_SIZE
)
(
    input clk, 
    input rst_n,
    input en,
    output done,
    input  [SIZE - 1:0] in0,
    input  [SIZE - 1:0] in1,
    input  [SIZE - 1:0] in2,
    input  [SIZE - 1:0] in3,
    input  [SIZE - 1:0] in4,
    input  [SIZE - 1:0] in5,
    input  [SIZE - 1:0] in6,
    input  [SIZE - 1:0] in7,
    input  [SIZE - 1:0] in8,
    input  [SIZE - 1:0] in9,
    input  [SIZE - 1:0] in10,
    input  [SIZE - 1:0] in11,
    input  [SIZE - 1:0] in12,
    input  [SIZE - 1:0] in13,
    input  [SIZE - 1:0] in14,
    input  [SIZE - 1:0] in15,
    input  [SIZE - 1:0] in16,
    input  [SIZE - 1:0] in17,
    input  [SIZE - 1:0] in18,
    input  [SIZE - 1:0] in19,
    input  [SIZE - 1:0] in20,
    input  [SIZE - 1:0] in21,
    input  [SIZE - 1:0] in22,
    input  [SIZE - 1:0] in23,
    input  [SIZE - 1:0] in24,
    input  [SIZE - 1:0] in25,
    input  [SIZE - 1:0] in26,
    input  [SIZE - 1:0] in27,
    input  [SIZE - 1:0] in28,
    input  [SIZE - 1:0] in29,
    input  [SIZE - 1:0] in30,
    input  [SIZE - 1:0] in31,
    input  [SIZE - 1:0] in32,
    input  [SIZE - 1:0] in33,
    input  [SIZE - 1:0] in34,
    input  [SIZE - 1:0] in35,
    input  [SIZE - 1:0] in36,
    input  [SIZE - 1:0] in37,
    input  [SIZE - 1:0] in38,
    input  [SIZE - 1:0] in39,
    input  [SIZE - 1:0] in40,
    input  [SIZE - 1:0] in41,
    input  [SIZE - 1:0] in42,
    input  [SIZE - 1:0] in43,
    input  [SIZE - 1:0] in44,
    input  [SIZE - 1:0] in45,
    input  [SIZE - 1:0] in46,
    input  [SIZE - 1:0] in47,
    input  [SIZE - 1:0] in48,
    input  [SIZE - 1:0] in49,
    input  [SIZE - 1:0] in50,
    input  [SIZE - 1:0] in51,
    input  [SIZE - 1:0] in52,
    input  [SIZE - 1:0] in53,
    input  [SIZE - 1:0] in54,
    input  [SIZE - 1:0] in55,
    input  [SIZE - 1:0] in56,
    input  [SIZE - 1:0] in57,
    input  [SIZE - 1:0] in58,
    input  [SIZE - 1:0] in59,
    input  [SIZE - 1:0] in60,
    input  [SIZE - 1:0] in61,
    input  [SIZE - 1:0] in62,
    input  [SIZE - 1:0] in63,
    input  [SIZE - 1:0] in64,
    input  [SIZE - 1:0] in65,
    input  [SIZE - 1:0] in66,
    input  [SIZE - 1:0] in67,
    input  [SIZE - 1:0] in68,
    input  [SIZE - 1:0] in69,
    input  [SIZE - 1:0] in70,
    input  [SIZE - 1:0] in71,
    input  [SIZE - 1:0] in72,
    input  [SIZE - 1:0] in73,
    input  [SIZE - 1:0] in74,
    input  [SIZE - 1:0] in75,
    input  [SIZE - 1:0] in76,
    input  [SIZE - 1:0] in77,
    input  [SIZE - 1:0] in78,
    input  [SIZE - 1:0] in79,
    input  [SIZE - 1:0] in80,
    input  [SIZE - 1:0] in81,
    input  [SIZE - 1:0] in82,
    input  [SIZE - 1:0] in83,
    input  [SIZE - 1:0] in84,
    input  [SIZE - 1:0] in85,
    input  [SIZE - 1:0] in86,
    input  [SIZE - 1:0] in87,
    input  [SIZE - 1:0] in88,
    input  [SIZE - 1:0] in89,
    input  [SIZE - 1:0] in90,
    input  [SIZE - 1:0] in91,
    input  [SIZE - 1:0] in92,
    input  [SIZE - 1:0] in93,
    input  [SIZE - 1:0] in94,
    input  [SIZE - 1:0] in95,
    input  [SIZE - 1:0] in96,
    input  [SIZE - 1:0] in97,
    input  [SIZE - 1:0] in98,
    input  [SIZE - 1:0] in99,
    input  [SIZE - 1:0] in100,
    input  [SIZE - 1:0] in101,
    input  [SIZE - 1:0] in102,
    input  [SIZE - 1:0] in103,
    input  [SIZE - 1:0] in104,
    input  [SIZE - 1:0] in105,
    input  [SIZE - 1:0] in106,
    input  [SIZE - 1:0] in107,
    input  [SIZE - 1:0] in108,
    input  [SIZE - 1:0] in109,
    input  [SIZE - 1:0] in110,
    input  [SIZE - 1:0] in111,
    input  [SIZE - 1:0] in112,
    input  [SIZE - 1:0] in113,
    input  [SIZE - 1:0] in114,
    input  [SIZE - 1:0] in115,
    input  [SIZE - 1:0] in116,
    input  [SIZE - 1:0] in117,
    input  [SIZE - 1:0] in118,
    input  [SIZE - 1:0] in119,
    input  [SIZE - 1:0] in120,
    input  [SIZE - 1:0] in121,
    input  [SIZE - 1:0] in122,
    input  [SIZE - 1:0] in123,
    input  [SIZE - 1:0] in124,
    input  [SIZE - 1:0] in125,
    input  [SIZE - 1:0] in126,
    input  [SIZE - 1:0] in127,
    input  [SIZE - 1:0] in128,
    input  [SIZE - 1:0] in129,
    input  [SIZE - 1:0] in130,
    input  [SIZE - 1:0] in131,
    input  [SIZE - 1:0] in132,
    input  [SIZE - 1:0] in133,
    input  [SIZE - 1:0] in134,
    input  [SIZE - 1:0] in135,
    input  [SIZE - 1:0] in136,
    input  [SIZE - 1:0] in137,
    input  [SIZE - 1:0] in138,
    input  [SIZE - 1:0] in139,
    input  [SIZE - 1:0] in140,
    input  [SIZE - 1:0] in141,
    input  [SIZE - 1:0] in142,
    input  [SIZE - 1:0] in143,
    input  [SIZE - 1:0] in144,
    input  [SIZE - 1:0] in145,
    input  [SIZE - 1:0] in146,
    input  [SIZE - 1:0] in147,
    input  [SIZE - 1:0] in148,
    input  [SIZE - 1:0] in149,
    input  [SIZE - 1:0] in150,
    input  [SIZE - 1:0] in151,
    input  [SIZE - 1:0] in152,
    input  [SIZE - 1:0] in153,
    input  [SIZE - 1:0] in154,
    input  [SIZE - 1:0] in155,
    input  [SIZE - 1:0] in156,
    input  [SIZE - 1:0] in157,
    input  [SIZE - 1:0] in158,
    input  [SIZE - 1:0] in159,
    input  [SIZE - 1:0] in160,
    input  [SIZE - 1:0] in161,
    input  [SIZE - 1:0] in162,
    input  [SIZE - 1:0] in163,
    input  [SIZE - 1:0] in164,
    input  [SIZE - 1:0] in165,
    input  [SIZE - 1:0] in166,
    input  [SIZE - 1:0] in167,
    input  [SIZE - 1:0] in168,
    input  [SIZE - 1:0] in169,
    input  [SIZE - 1:0] in170,
    input  [SIZE - 1:0] in171,
    input  [SIZE - 1:0] in172,
    input  [SIZE - 1:0] in173,
    input  [SIZE - 1:0] in174,
    input  [SIZE - 1:0] in175,
    input  [SIZE - 1:0] in176,
    input  [SIZE - 1:0] in177,
    input  [SIZE - 1:0] in178,
    input  [SIZE - 1:0] in179,
    input  [SIZE - 1:0] in180,
    input  [SIZE - 1:0] in181,
    input  [SIZE - 1:0] in182,
    input  [SIZE - 1:0] in183,
    input  [SIZE - 1:0] in184,
    input  [SIZE - 1:0] in185,
    input  [SIZE - 1:0] in186,
    input  [SIZE - 1:0] in187,
    input  [SIZE - 1:0] in188,
    input  [SIZE - 1:0] in189,
    input  [SIZE - 1:0] in190,
    input  [SIZE - 1:0] in191,
    input  [SIZE - 1:0] in192,
    input  [SIZE - 1:0] in193,
    input  [SIZE - 1:0] in194,
    input  [SIZE - 1:0] in195,
    input  [SIZE - 1:0] in196,
    input  [SIZE - 1:0] in197,
    input  [SIZE - 1:0] in198,
    input  [SIZE - 1:0] in199,
    input  [SIZE - 1:0] in200,
    input  [SIZE - 1:0] in201,
    input  [SIZE - 1:0] in202,
    input  [SIZE - 1:0] in203,
    input  [SIZE - 1:0] in204,
    input  [SIZE - 1:0] in205,
    input  [SIZE - 1:0] in206,
    input  [SIZE - 1:0] in207,
    input  [SIZE - 1:0] in208,
    input  [SIZE - 1:0] in209,
    input  [SIZE - 1:0] in210,
    input  [SIZE - 1:0] in211,
    input  [SIZE - 1:0] in212,
    input  [SIZE - 1:0] in213,
    input  [SIZE - 1:0] in214,
    input  [SIZE - 1:0] in215,
    input  [SIZE - 1:0] in216,
    input  [SIZE - 1:0] in217,
    input  [SIZE - 1:0] in218,
    input  [SIZE - 1:0] in219,
    input  [SIZE - 1:0] in220,
    input  [SIZE - 1:0] in221,
    input  [SIZE - 1:0] in222,
    input  [SIZE - 1:0] in223,
    input  [SIZE - 1:0] in224,
    input  [SIZE - 1:0] in225,
    input  [SIZE - 1:0] in226,
    input  [SIZE - 1:0] in227,
    input  [SIZE - 1:0] in228,
    input  [SIZE - 1:0] in229,
    input  [SIZE - 1:0] in230,
    input  [SIZE - 1:0] in231,
    input  [SIZE - 1:0] in232,
    input  [SIZE - 1:0] in233,
    input  [SIZE - 1:0] in234,
    input  [SIZE - 1:0] in235,
    input  [SIZE - 1:0] in236,
    input  [SIZE - 1:0] in237,
    input  [SIZE - 1:0] in238,
    input  [SIZE - 1:0] in239,
    input  [SIZE - 1:0] in240,
    input  [SIZE - 1:0] in241,
    input  [SIZE - 1:0] in242,
    input  [SIZE - 1:0] in243,
    input  [SIZE - 1:0] in244,
    input  [SIZE - 1:0] in245,
    input  [SIZE - 1:0] in246,
    input  [SIZE - 1:0] in247,
    input  [SIZE - 1:0] in248,
    input  [SIZE - 1:0] in249,
    input  [SIZE - 1:0] in250,
    input  [SIZE - 1:0] in251,
    input  [SIZE - 1:0] in252,
    input  [SIZE - 1:0] in253,
    input  [SIZE - 1:0] in254,
    input  [SIZE - 1:0] in255,
    input  [SIZE - 1:0] in256,
    input  [SIZE - 1:0] in257,
    input  [SIZE - 1:0] in258,
    input  [SIZE - 1:0] in259,
    input  [SIZE - 1:0] in260,
    input  [SIZE - 1:0] in261,
    input  [SIZE - 1:0] in262,
    input  [SIZE - 1:0] in263,
    input  [SIZE - 1:0] in264,
    input  [SIZE - 1:0] in265,
    input  [SIZE - 1:0] in266,
    input  [SIZE - 1:0] in267,
    input  [SIZE - 1:0] in268,
    input  [SIZE - 1:0] in269,
    input  [SIZE - 1:0] in270,
    input  [SIZE - 1:0] in271,
    input  [SIZE - 1:0] in272,
    input  [SIZE - 1:0] in273,
    input  [SIZE - 1:0] in274,
    input  [SIZE - 1:0] in275,
    input  [SIZE - 1:0] in276,
    input  [SIZE - 1:0] in277,
    input  [SIZE - 1:0] in278,
    input  [SIZE - 1:0] in279,
    input  [SIZE - 1:0] in280,
    input  [SIZE - 1:0] in281,
    input  [SIZE - 1:0] in282,
    input  [SIZE - 1:0] in283,
    input  [SIZE - 1:0] in284,
    input  [SIZE - 1:0] in285,
    input  [SIZE - 1:0] in286,
    input  [SIZE - 1:0] in287,
    input  [SIZE - 1:0] in288,
    input  [SIZE - 1:0] in289,
    input  [SIZE - 1:0] in290,
    input  [SIZE - 1:0] in291,
    input  [SIZE - 1:0] in292,
    input  [SIZE - 1:0] in293,
    input  [SIZE - 1:0] in294,
    input  [SIZE - 1:0] in295,
    input  [SIZE - 1:0] in296,
    input  [SIZE - 1:0] in297,
    input  [SIZE - 1:0] in298,
    input  [SIZE - 1:0] in299,
    input  [SIZE - 1:0] in300,
    input  [SIZE - 1:0] in301,
    input  [SIZE - 1:0] in302,
    input  [SIZE - 1:0] in303,
    input  [SIZE - 1:0] in304,
    input  [SIZE - 1:0] in305,
    input  [SIZE - 1:0] in306,
    input  [SIZE - 1:0] in307,
    input  [SIZE - 1:0] in308,
    input  [SIZE - 1:0] in309,
    input  [SIZE - 1:0] in310,
    input  [SIZE - 1:0] in311,
    input  [SIZE - 1:0] in312,
    input  [SIZE - 1:0] in313,
    input  [SIZE - 1:0] in314,
    input  [SIZE - 1:0] in315,
    input  [SIZE - 1:0] in316,
    input  [SIZE - 1:0] in317,
    input  [SIZE - 1:0] in318,
    input  [SIZE - 1:0] in319,
    input  [SIZE - 1:0] in320,
    input  [SIZE - 1:0] in321,
    input  [SIZE - 1:0] in322,
    input  [SIZE - 1:0] in323,
    input  [SIZE - 1:0] in324,
    input  [SIZE - 1:0] in325,
    input  [SIZE - 1:0] in326,
    input  [SIZE - 1:0] in327,
    input  [SIZE - 1:0] in328,
    input  [SIZE - 1:0] in329,
    input  [SIZE - 1:0] in330,
    input  [SIZE - 1:0] in331,
    input  [SIZE - 1:0] in332,
    input  [SIZE - 1:0] in333,
    input  [SIZE - 1:0] in334,
    input  [SIZE - 1:0] in335,
    input  [SIZE - 1:0] in336,
    input  [SIZE - 1:0] in337,
    input  [SIZE - 1:0] in338,
    input  [SIZE - 1:0] in339,
    input  [SIZE - 1:0] in340,
    input  [SIZE - 1:0] in341,
    input  [SIZE - 1:0] in342,
    input  [SIZE - 1:0] in343,
    input  [SIZE - 1:0] in344,
    input  [SIZE - 1:0] in345,
    input  [SIZE - 1:0] in346,
    input  [SIZE - 1:0] in347,
    input  [SIZE - 1:0] in348,
    input  [SIZE - 1:0] in349,
    input  [SIZE - 1:0] in350,
    input  [SIZE - 1:0] in351,
    input  [SIZE - 1:0] in352,
    input  [SIZE - 1:0] in353,
    input  [SIZE - 1:0] in354,
    input  [SIZE - 1:0] in355,
    input  [SIZE - 1:0] in356,
    input  [SIZE - 1:0] in357,
    input  [SIZE - 1:0] in358,
    input  [SIZE - 1:0] in359,
    input  [SIZE - 1:0] in360,
    input  [SIZE - 1:0] in361,
    input  [SIZE - 1:0] in362,
    input  [SIZE - 1:0] in363,
    input  [SIZE - 1:0] in364,
    input  [SIZE - 1:0] in365,
    input  [SIZE - 1:0] in366,
    input  [SIZE - 1:0] in367,
    input  [SIZE - 1:0] in368,
    input  [SIZE - 1:0] in369,
    input  [SIZE - 1:0] in370,
    input  [SIZE - 1:0] in371,
    input  [SIZE - 1:0] in372,
    input  [SIZE - 1:0] in373,
    input  [SIZE - 1:0] in374,
    input  [SIZE - 1:0] in375,
    input  [SIZE - 1:0] in376,
    input  [SIZE - 1:0] in377,
    input  [SIZE - 1:0] in378,
    input  [SIZE - 1:0] in379,
    input  [SIZE - 1:0] in380,
    input  [SIZE - 1:0] in381,
    input  [SIZE - 1:0] in382,
    input  [SIZE - 1:0] in383,
    input  [SIZE - 1:0] in384,
    input  [SIZE - 1:0] in385,
    input  [SIZE - 1:0] in386,
    input  [SIZE - 1:0] in387,
    input  [SIZE - 1:0] in388,
    input  [SIZE - 1:0] in389,
    input  [SIZE - 1:0] in390,
    input  [SIZE - 1:0] in391,
    input  [SIZE - 1:0] in392,
    input  [SIZE - 1:0] in393,
    input  [SIZE - 1:0] in394,
    input  [SIZE - 1:0] in395,
    input  [SIZE - 1:0] in396,
    input  [SIZE - 1:0] in397,
    input  [SIZE - 1:0] in398,
    input  [SIZE - 1:0] in399,
    input  [SIZE - 1:0] in400,
    input  [SIZE - 1:0] in401,
    input  [SIZE - 1:0] in402,
    input  [SIZE - 1:0] in403,
    input  [SIZE - 1:0] in404,
    input  [SIZE - 1:0] in405,
    input  [SIZE - 1:0] in406,
    input  [SIZE - 1:0] in407,
    input  [SIZE - 1:0] in408,
    input  [SIZE - 1:0] in409,
    input  [SIZE - 1:0] in410,
    input  [SIZE - 1:0] in411,
    input  [SIZE - 1:0] in412,
    input  [SIZE - 1:0] in413,
    input  [SIZE - 1:0] in414,
    input  [SIZE - 1:0] in415,
    input  [SIZE - 1:0] in416,
    input  [SIZE - 1:0] in417,
    input  [SIZE - 1:0] in418,
    input  [SIZE - 1:0] in419,
    input  [SIZE - 1:0] in420,
    input  [SIZE - 1:0] in421,
    input  [SIZE - 1:0] in422,
    input  [SIZE - 1:0] in423,
    input  [SIZE - 1:0] in424,
    input  [SIZE - 1:0] in425,
    input  [SIZE - 1:0] in426,
    input  [SIZE - 1:0] in427,
    input  [SIZE - 1:0] in428,
    input  [SIZE - 1:0] in429,
    input  [SIZE - 1:0] in430,
    input  [SIZE - 1:0] in431,
    input  [SIZE - 1:0] in432,
    input  [SIZE - 1:0] in433,
    input  [SIZE - 1:0] in434,
    input  [SIZE - 1:0] in435,
    input  [SIZE - 1:0] in436,
    input  [SIZE - 1:0] in437,
    input  [SIZE - 1:0] in438,
    input  [SIZE - 1:0] in439,
    input  [SIZE - 1:0] in440,
    input  [SIZE - 1:0] in441,
    input  [SIZE - 1:0] in442,
    input  [SIZE - 1:0] in443,
    input  [SIZE - 1:0] in444,
    input  [SIZE - 1:0] in445,
    input  [SIZE - 1:0] in446,
    input  [SIZE - 1:0] in447,
    input  [SIZE - 1:0] in448,
    input  [SIZE - 1:0] in449,
    input  [SIZE - 1:0] in450,
    input  [SIZE - 1:0] in451,
    input  [SIZE - 1:0] in452,
    input  [SIZE - 1:0] in453,
    input  [SIZE - 1:0] in454,
    input  [SIZE - 1:0] in455,
    input  [SIZE - 1:0] in456,
    input  [SIZE - 1:0] in457,
    input  [SIZE - 1:0] in458,
    input  [SIZE - 1:0] in459,
    input  [SIZE - 1:0] in460,
    input  [SIZE - 1:0] in461,
    input  [SIZE - 1:0] in462,
    input  [SIZE - 1:0] in463,
    input  [SIZE - 1:0] in464,
    input  [SIZE - 1:0] in465,
    input  [SIZE - 1:0] in466,
    input  [SIZE - 1:0] in467,
    input  [SIZE - 1:0] in468,
    input  [SIZE - 1:0] in469,
    input  [SIZE - 1:0] in470,
    input  [SIZE - 1:0] in471,
    input  [SIZE - 1:0] in472,
    input  [SIZE - 1:0] in473,
    input  [SIZE - 1:0] in474,
    input  [SIZE - 1:0] in475,
    input  [SIZE - 1:0] in476,
    input  [SIZE - 1:0] in477,
    input  [SIZE - 1:0] in478,
    input  [SIZE - 1:0] in479,
    input  [SIZE - 1:0] in480,
    input  [SIZE - 1:0] in481,
    input  [SIZE - 1:0] in482,
    input  [SIZE - 1:0] in483,
    input  [SIZE - 1:0] in484,
    input  [SIZE - 1:0] in485,
    input  [SIZE - 1:0] in486,
    input  [SIZE - 1:0] in487,
    input  [SIZE - 1:0] in488,
    input  [SIZE - 1:0] in489,
    input  [SIZE - 1:0] in490,
    input  [SIZE - 1:0] in491,
    input  [SIZE - 1:0] in492,
    input  [SIZE - 1:0] in493,
    input  [SIZE - 1:0] in494,
    input  [SIZE - 1:0] in495,
    input  [SIZE - 1:0] in496,
    input  [SIZE - 1:0] in497,
    input  [SIZE - 1:0] in498,
    input  [SIZE - 1:0] in499,
    input  [SIZE - 1:0] in500,
    input  [SIZE - 1:0] in501,
    input  [SIZE - 1:0] in502,
    input  [SIZE - 1:0] in503,
    input  [SIZE - 1:0] in504,
    input  [SIZE - 1:0] in505,
    input  [SIZE - 1:0] in506,
    input  [SIZE - 1:0] in507,
    input  [SIZE - 1:0] in508,
    input  [SIZE - 1:0] in509,
    input  [SIZE - 1:0] in510,
    input  [SIZE - 1:0] in511,
    input  [SIZE - 1:0] in512,
    input  [SIZE - 1:0] in513,
    input  [SIZE - 1:0] in514,
    input  [SIZE - 1:0] in515,
    input  [SIZE - 1:0] in516,
    input  [SIZE - 1:0] in517,
    input  [SIZE - 1:0] in518,
    input  [SIZE - 1:0] in519,
    input  [SIZE - 1:0] in520,
    input  [SIZE - 1:0] in521,
    input  [SIZE - 1:0] in522,
    input  [SIZE - 1:0] in523,
    input  [SIZE - 1:0] in524,
    input  [SIZE - 1:0] in525,
    input  [SIZE - 1:0] in526,
    input  [SIZE - 1:0] in527,
    input  [SIZE - 1:0] in528,
    input  [SIZE - 1:0] in529,
    input  [SIZE - 1:0] in530,
    input  [SIZE - 1:0] in531,
    input  [SIZE - 1:0] in532,
    input  [SIZE - 1:0] in533,
    input  [SIZE - 1:0] in534,
    input  [SIZE - 1:0] in535,
    input  [SIZE - 1:0] in536,
    input  [SIZE - 1:0] in537,
    input  [SIZE - 1:0] in538,
    input  [SIZE - 1:0] in539,
    input  [SIZE - 1:0] in540,
    input  [SIZE - 1:0] in541,
    input  [SIZE - 1:0] in542,
    input  [SIZE - 1:0] in543,
    input  [SIZE - 1:0] in544,
    input  [SIZE - 1:0] in545,
    input  [SIZE - 1:0] in546,
    input  [SIZE - 1:0] in547,
    input  [SIZE - 1:0] in548,
    input  [SIZE - 1:0] in549,
    input  [SIZE - 1:0] in550,
    input  [SIZE - 1:0] in551,
    input  [SIZE - 1:0] in552,
    input  [SIZE - 1:0] in553,
    input  [SIZE - 1:0] in554,
    input  [SIZE - 1:0] in555,
    input  [SIZE - 1:0] in556,
    input  [SIZE - 1:0] in557,
    input  [SIZE - 1:0] in558,
    input  [SIZE - 1:0] in559,
    input  [SIZE - 1:0] in560,
    input  [SIZE - 1:0] in561,
    input  [SIZE - 1:0] in562,
    input  [SIZE - 1:0] in563,
    input  [SIZE - 1:0] in564,
    input  [SIZE - 1:0] in565,
    input  [SIZE - 1:0] in566,
    input  [SIZE - 1:0] in567,
    input  [SIZE - 1:0] in568,
    input  [SIZE - 1:0] in569,
    input  [SIZE - 1:0] in570,
    input  [SIZE - 1:0] in571,
    input  [SIZE - 1:0] in572,
    input  [SIZE - 1:0] in573,
    input  [SIZE - 1:0] in574,
    input  [SIZE - 1:0] in575,
    input  [SIZE - 1:0] in576,
    input  [SIZE - 1:0] in577,
    input  [SIZE - 1:0] in578,
    input  [SIZE - 1:0] in579,
    input  [SIZE - 1:0] in580,
    input  [SIZE - 1:0] in581,
    input  [SIZE - 1:0] in582,
    input  [SIZE - 1:0] in583,
    input  [SIZE - 1:0] in584,
    input  [SIZE - 1:0] in585,
    input  [SIZE - 1:0] in586,
    input  [SIZE - 1:0] in587,
    input  [SIZE - 1:0] in588,
    input  [SIZE - 1:0] in589,
    input  [SIZE - 1:0] in590,
    input  [SIZE - 1:0] in591,
    input  [SIZE - 1:0] in592,
    input  [SIZE - 1:0] in593,
    input  [SIZE - 1:0] in594,
    input  [SIZE - 1:0] in595,
    input  [SIZE - 1:0] in596,
    input  [SIZE - 1:0] in597,
    input  [SIZE - 1:0] in598,
    input  [SIZE - 1:0] in599,
    input  [SIZE - 1:0] in600,
    input  [SIZE - 1:0] in601,
    input  [SIZE - 1:0] in602,
    input  [SIZE - 1:0] in603,
    input  [SIZE - 1:0] in604,
    input  [SIZE - 1:0] in605,
    input  [SIZE - 1:0] in606,
    input  [SIZE - 1:0] in607,
    input  [SIZE - 1:0] in608,
    input  [SIZE - 1:0] in609,
    input  [SIZE - 1:0] in610,
    input  [SIZE - 1:0] in611,
    input  [SIZE - 1:0] in612,
    input  [SIZE - 1:0] in613,
    input  [SIZE - 1:0] in614,
    input  [SIZE - 1:0] in615,
    input  [SIZE - 1:0] in616,
    input  [SIZE - 1:0] in617,
    input  [SIZE - 1:0] in618,
    input  [SIZE - 1:0] in619,
    input  [SIZE - 1:0] in620,
    input  [SIZE - 1:0] in621,
    input  [SIZE - 1:0] in622,
    input  [SIZE - 1:0] in623,
    input  [SIZE - 1:0] in624,
    input  [SIZE - 1:0] in625,
    input  [SIZE - 1:0] in626,
    input  [SIZE - 1:0] in627,
    input  [SIZE - 1:0] in628,
    input  [SIZE - 1:0] in629,
    input  [SIZE - 1:0] in630,
    input  [SIZE - 1:0] in631,
    input  [SIZE - 1:0] in632,
    input  [SIZE - 1:0] in633,
    input  [SIZE - 1:0] in634,
    input  [SIZE - 1:0] in635,
    input  [SIZE - 1:0] in636,
    input  [SIZE - 1:0] in637,
    input  [SIZE - 1:0] in638,
    input  [SIZE - 1:0] in639,
    input  [SIZE - 1:0] in640,
    input  [SIZE - 1:0] in641,
    input  [SIZE - 1:0] in642,
    input  [SIZE - 1:0] in643,
    input  [SIZE - 1:0] in644,
    input  [SIZE - 1:0] in645,
    input  [SIZE - 1:0] in646,
    input  [SIZE - 1:0] in647,
    input  [SIZE - 1:0] in648,
    input  [SIZE - 1:0] in649,
    input  [SIZE - 1:0] in650,
    input  [SIZE - 1:0] in651,
    input  [SIZE - 1:0] in652,
    input  [SIZE - 1:0] in653,
    input  [SIZE - 1:0] in654,
    input  [SIZE - 1:0] in655,
    input  [SIZE - 1:0] in656,
    input  [SIZE - 1:0] in657,
    input  [SIZE - 1:0] in658,
    input  [SIZE - 1:0] in659,
    input  [SIZE - 1:0] in660,
    input  [SIZE - 1:0] in661,
    input  [SIZE - 1:0] in662,
    input  [SIZE - 1:0] in663,
    input  [SIZE - 1:0] in664,
    input  [SIZE - 1:0] in665,
    input  [SIZE - 1:0] in666,
    input  [SIZE - 1:0] in667,
    input  [SIZE - 1:0] in668,
    input  [SIZE - 1:0] in669,
    input  [SIZE - 1:0] in670,
    input  [SIZE - 1:0] in671,
    input  [SIZE - 1:0] in672,
    input  [SIZE - 1:0] in673,
    input  [SIZE - 1:0] in674,
    input  [SIZE - 1:0] in675,
    input  [SIZE - 1:0] in676,
    input  [SIZE - 1:0] in677,
    input  [SIZE - 1:0] in678,
    input  [SIZE - 1:0] in679,
    input  [SIZE - 1:0] in680,
    input  [SIZE - 1:0] in681,
    input  [SIZE - 1:0] in682,
    input  [SIZE - 1:0] in683,
    input  [SIZE - 1:0] in684,
    input  [SIZE - 1:0] in685,
    input  [SIZE - 1:0] in686,
    input  [SIZE - 1:0] in687,
    input  [SIZE - 1:0] in688,
    input  [SIZE - 1:0] in689,
    input  [SIZE - 1:0] in690,
    input  [SIZE - 1:0] in691,
    input  [SIZE - 1:0] in692,
    input  [SIZE - 1:0] in693,
    input  [SIZE - 1:0] in694,
    input  [SIZE - 1:0] in695,
    input  [SIZE - 1:0] in696,
    input  [SIZE - 1:0] in697,
    input  [SIZE - 1:0] in698,
    input  [SIZE - 1:0] in699,
    input  [SIZE - 1:0] in700,
    input  [SIZE - 1:0] in701,
    input  [SIZE - 1:0] in702,
    input  [SIZE - 1:0] in703,
    input  [SIZE - 1:0] in704,
    input  [SIZE - 1:0] in705,
    input  [SIZE - 1:0] in706,
    input  [SIZE - 1:0] in707,
    input  [SIZE - 1:0] in708,
    input  [SIZE - 1:0] in709,
    input  [SIZE - 1:0] in710,
    input  [SIZE - 1:0] in711,
    input  [SIZE - 1:0] in712,
    input  [SIZE - 1:0] in713,
    input  [SIZE - 1:0] in714,
    input  [SIZE - 1:0] in715,
    input  [SIZE - 1:0] in716,
    input  [SIZE - 1:0] in717,
    input  [SIZE - 1:0] in718,
    input  [SIZE - 1:0] in719,
    input  [SIZE - 1:0] in720,
    input  [SIZE - 1:0] in721,
    input  [SIZE - 1:0] in722,
    input  [SIZE - 1:0] in723,
    input  [SIZE - 1:0] in724,
    input  [SIZE - 1:0] in725,
    input  [SIZE - 1:0] in726,
    input  [SIZE - 1:0] in727,
    input  [SIZE - 1:0] in728,
    input  [SIZE - 1:0] in729,
    input  [SIZE - 1:0] in730,
    input  [SIZE - 1:0] in731,
    input  [SIZE - 1:0] in732,
    input  [SIZE - 1:0] in733,
    input  [SIZE - 1:0] in734,
    input  [SIZE - 1:0] in735,
    input  [SIZE - 1:0] in736,
    input  [SIZE - 1:0] in737,
    input  [SIZE - 1:0] in738,
    input  [SIZE - 1:0] in739,
    input  [SIZE - 1:0] in740,
    input  [SIZE - 1:0] in741,
    input  [SIZE - 1:0] in742,
    input  [SIZE - 1:0] in743,
    input  [SIZE - 1:0] in744,
    input  [SIZE - 1:0] in745,
    input  [SIZE - 1:0] in746,
    input  [SIZE - 1:0] in747,
    input  [SIZE - 1:0] in748,
    input  [SIZE - 1:0] in749,
    input  [SIZE - 1:0] in750,
    input  [SIZE - 1:0] in751,
    input  [SIZE - 1:0] in752,
    input  [SIZE - 1:0] in753,
    input  [SIZE - 1:0] in754,
    input  [SIZE - 1:0] in755,
    input  [SIZE - 1:0] in756,
    input  [SIZE - 1:0] in757,
    input  [SIZE - 1:0] in758,
    input  [SIZE - 1:0] in759,
    input  [SIZE - 1:0] in760,
    input  [SIZE - 1:0] in761,
    input  [SIZE - 1:0] in762,
    input  [SIZE - 1:0] in763,
    input  [SIZE - 1:0] in764,
    input  [SIZE - 1:0] in765,
    input  [SIZE - 1:0] in766,
    input  [SIZE - 1:0] in767,
    input  [SIZE - 1:0] in768,
    input  [SIZE - 1:0] in769,
    input  [SIZE - 1:0] in770,
    input  [SIZE - 1:0] in771,
    input  [SIZE - 1:0] in772,
    input  [SIZE - 1:0] in773,
    input  [SIZE - 1:0] in774,
    input  [SIZE - 1:0] in775,
    input  [SIZE - 1:0] in776,
    input  [SIZE - 1:0] in777,
    input  [SIZE - 1:0] in778,
    input  [SIZE - 1:0] in779,
    input  [SIZE - 1:0] in780,
    input  [SIZE - 1:0] in781,
    input  [SIZE - 1:0] in782,
    input  [SIZE - 1:0] in783,
    input  [SIZE - 1:0] in784,
    input  [SIZE - 1:0] in785,
    input  [SIZE - 1:0] in786,
    input  [SIZE - 1:0] in787,
    input  [SIZE - 1:0] in788,
    input  [SIZE - 1:0] in789,
    input  [SIZE - 1:0] in790,
    input  [SIZE - 1:0] in791,
    input  [SIZE - 1:0] in792,
    input  [SIZE - 1:0] in793,
    input  [SIZE - 1:0] in794,
    input  [SIZE - 1:0] in795,
    input  [SIZE - 1:0] in796,
    input  [SIZE - 1:0] in797,
    input  [SIZE - 1:0] in798,
    input  [SIZE - 1:0] in799,
    input  [SIZE - 1:0] in800,
    input  [SIZE - 1:0] in801,
    input  [SIZE - 1:0] in802,
    input  [SIZE - 1:0] in803,
    input  [SIZE - 1:0] in804,
    input  [SIZE - 1:0] in805,
    input  [SIZE - 1:0] in806,
    input  [SIZE - 1:0] in807,
    input  [SIZE - 1:0] in808,
    input  [SIZE - 1:0] in809,
    input  [SIZE - 1:0] in810,
    input  [SIZE - 1:0] in811,
    input  [SIZE - 1:0] in812,
    input  [SIZE - 1:0] in813,
    input  [SIZE - 1:0] in814,
    input  [SIZE - 1:0] in815,
    input  [SIZE - 1:0] in816,
    input  [SIZE - 1:0] in817,
    input  [SIZE - 1:0] in818,
    input  [SIZE - 1:0] in819,
    input  [SIZE - 1:0] in820,
    input  [SIZE - 1:0] in821,
    input  [SIZE - 1:0] in822,
    input  [SIZE - 1:0] in823,
    input  [SIZE - 1:0] in824,
    input  [SIZE - 1:0] in825,
    input  [SIZE - 1:0] in826,
    input  [SIZE - 1:0] in827,
    input  [SIZE - 1:0] in828,
    input  [SIZE - 1:0] in829,
    input  [SIZE - 1:0] in830,
    input  [SIZE - 1:0] in831,
    input  [SIZE - 1:0] in832,
    input  [SIZE - 1:0] in833,
    input  [SIZE - 1:0] in834,
    input  [SIZE - 1:0] in835,
    input  [SIZE - 1:0] in836,
    input  [SIZE - 1:0] in837,
    input  [SIZE - 1:0] in838,
    input  [SIZE - 1:0] in839,
    input  [SIZE - 1:0] in840,
    input  [SIZE - 1:0] in841,
    input  [SIZE - 1:0] in842,
    input  [SIZE - 1:0] in843,
    input  [SIZE - 1:0] in844,
    input  [SIZE - 1:0] in845,
    input  [SIZE - 1:0] in846,
    input  [SIZE - 1:0] in847,
    input  [SIZE - 1:0] in848,
    input  [SIZE - 1:0] in849,
    input  [SIZE - 1:0] in850,
    input  [SIZE - 1:0] in851,
    input  [SIZE - 1:0] in852,
    input  [SIZE - 1:0] in853,
    input  [SIZE - 1:0] in854,
    input  [SIZE - 1:0] in855,
    input  [SIZE - 1:0] in856,
    input  [SIZE - 1:0] in857,
    input  [SIZE - 1:0] in858,
    input  [SIZE - 1:0] in859,
    input  [SIZE - 1:0] in860,
    input  [SIZE - 1:0] in861,
    input  [SIZE - 1:0] in862,
    input  [SIZE - 1:0] in863,
    input  [SIZE - 1:0] in864,
    input  [SIZE - 1:0] in865,
    input  [SIZE - 1:0] in866,
    input  [SIZE - 1:0] in867,
    input  [SIZE - 1:0] in868,
    input  [SIZE - 1:0] in869,
    input  [SIZE - 1:0] in870,
    input  [SIZE - 1:0] in871,
    input  [SIZE - 1:0] in872,
    input  [SIZE - 1:0] in873,
    input  [SIZE - 1:0] in874,
    input  [SIZE - 1:0] in875,
    input  [SIZE - 1:0] in876,
    input  [SIZE - 1:0] in877,
    input  [SIZE - 1:0] in878,
    input  [SIZE - 1:0] in879,
    input  [SIZE - 1:0] in880,
    input  [SIZE - 1:0] in881,
    input  [SIZE - 1:0] in882,
    input  [SIZE - 1:0] in883,
    input  [SIZE - 1:0] in884,
    input  [SIZE - 1:0] in885,
    input  [SIZE - 1:0] in886,
    input  [SIZE - 1:0] in887,
    input  [SIZE - 1:0] in888,
    input  [SIZE - 1:0] in889,
    input  [SIZE - 1:0] in890,
    input  [SIZE - 1:0] in891,
    input  [SIZE - 1:0] in892,
    input  [SIZE - 1:0] in893,
    input  [SIZE - 1:0] in894,
    input  [SIZE - 1:0] in895,
    input  [SIZE - 1:0] in896,
    input  [SIZE - 1:0] in897,
    input  [SIZE - 1:0] in898,
    input  [SIZE - 1:0] in899,
    input  [SIZE - 1:0] in900,
    input  [SIZE - 1:0] in901,
    input  [SIZE - 1:0] in902,
    input  [SIZE - 1:0] in903,
    input  [SIZE - 1:0] in904,
    input  [SIZE - 1:0] in905,
    input  [SIZE - 1:0] in906,
    input  [SIZE - 1:0] in907,
    input  [SIZE - 1:0] in908,
    input  [SIZE - 1:0] in909,
    input  [SIZE - 1:0] in910,
    input  [SIZE - 1:0] in911,
    input  [SIZE - 1:0] in912,
    input  [SIZE - 1:0] in913,
    input  [SIZE - 1:0] in914,
    input  [SIZE - 1:0] in915,
    input  [SIZE - 1:0] in916,
    input  [SIZE - 1:0] in917,
    input  [SIZE - 1:0] in918,
    input  [SIZE - 1:0] in919,
    input  [SIZE - 1:0] in920,
    input  [SIZE - 1:0] in921,
    input  [SIZE - 1:0] in922,
    input  [SIZE - 1:0] in923,
    input  [SIZE - 1:0] in924,
    input  [SIZE - 1:0] in925,
    input  [SIZE - 1:0] in926,
    input  [SIZE - 1:0] in927,
    input  [SIZE - 1:0] in928,
    input  [SIZE - 1:0] in929,
    input  [SIZE - 1:0] in930,
    input  [SIZE - 1:0] in931,
    input  [SIZE - 1:0] in932,
    input  [SIZE - 1:0] in933,
    input  [SIZE - 1:0] in934,
    input  [SIZE - 1:0] in935,
    input  [SIZE - 1:0] in936,
    input  [SIZE - 1:0] in937,
    input  [SIZE - 1:0] in938,
    input  [SIZE - 1:0] in939,
    input  [SIZE - 1:0] in940,
    input  [SIZE - 1:0] in941,
    input  [SIZE - 1:0] in942,
    input  [SIZE - 1:0] in943,
    input  [SIZE - 1:0] in944,
    input  [SIZE - 1:0] in945,
    input  [SIZE - 1:0] in946,
    input  [SIZE - 1:0] in947,
    input  [SIZE - 1:0] in948,
    input  [SIZE - 1:0] in949,
    input  [SIZE - 1:0] in950,
    input  [SIZE - 1:0] in951,
    input  [SIZE - 1:0] in952,
    input  [SIZE - 1:0] in953,
    input  [SIZE - 1:0] in954,
    input  [SIZE - 1:0] in955,
    input  [SIZE - 1:0] in956,
    input  [SIZE - 1:0] in957,
    input  [SIZE - 1:0] in958,
    input  [SIZE - 1:0] in959,
    input  [SIZE - 1:0] in960,
    input  [SIZE - 1:0] in961,
    input  [SIZE - 1:0] in962,
    input  [SIZE - 1:0] in963,
    input  [SIZE - 1:0] in964,
    input  [SIZE - 1:0] in965,
    input  [SIZE - 1:0] in966,
    input  [SIZE - 1:0] in967,
    input  [SIZE - 1:0] in968,
    input  [SIZE - 1:0] in969,
    input  [SIZE - 1:0] in970,
    input  [SIZE - 1:0] in971,
    input  [SIZE - 1:0] in972,
    input  [SIZE - 1:0] in973,
    input  [SIZE - 1:0] in974,
    input  [SIZE - 1:0] in975,
    input  [SIZE - 1:0] in976,
    input  [SIZE - 1:0] in977,
    input  [SIZE - 1:0] in978,
    input  [SIZE - 1:0] in979,
    input  [SIZE - 1:0] in980,
    input  [SIZE - 1:0] in981,
    input  [SIZE - 1:0] in982,
    input  [SIZE - 1:0] in983,
    input  [SIZE - 1:0] in984,
    input  [SIZE - 1:0] in985,
    input  [SIZE - 1:0] in986,
    input  [SIZE - 1:0] in987,
    input  [SIZE - 1:0] in988,
    input  [SIZE - 1:0] in989,
    input  [SIZE - 1:0] in990,
    input  [SIZE - 1:0] in991,
    input  [SIZE - 1:0] in992,
    input  [SIZE - 1:0] in993,
    input  [SIZE - 1:0] in994,
    input  [SIZE - 1:0] in995,
    input  [SIZE - 1:0] in996,
    input  [SIZE - 1:0] in997,
    input  [SIZE - 1:0] in998,
    input  [SIZE - 1:0] in999,
    input  [SIZE - 1:0] in1000,
    input  [SIZE - 1:0] in1001,
    input  [SIZE - 1:0] in1002,
    input  [SIZE - 1:0] in1003,
    input  [SIZE - 1:0] in1004,
    input  [SIZE - 1:0] in1005,
    input  [SIZE - 1:0] in1006,
    input  [SIZE - 1:0] in1007,
    input  [SIZE - 1:0] in1008,
    input  [SIZE - 1:0] in1009,
    input  [SIZE - 1:0] in1010,
    input  [SIZE - 1:0] in1011,
    input  [SIZE - 1:0] in1012,
    input  [SIZE - 1:0] in1013,
    input  [SIZE - 1:0] in1014,
    input  [SIZE - 1:0] in1015,
    input  [SIZE - 1:0] in1016,
    input  [SIZE - 1:0] in1017,
    input  [SIZE - 1:0] in1018,
    input  [SIZE - 1:0] in1019,
    input  [SIZE - 1:0] in1020,
    input  [SIZE - 1:0] in1021,
    input  [SIZE - 1:0] in1022,
    input  [SIZE - 1:0] in1023,

    output [SIZE - 1:0] out0,
    output [SIZE - 1:0] out1,
    output [SIZE - 1:0] out2,
    output [SIZE - 1:0] out3,
    output [SIZE - 1:0] out4,
    output [SIZE - 1:0] out5,
    output [SIZE - 1:0] out6,
    output [SIZE - 1:0] out7,
    output [SIZE - 1:0] out8,
    output [SIZE - 1:0] out9,
    output [SIZE - 1:0] out10,
    output [SIZE - 1:0] out11,
    output [SIZE - 1:0] out12,
    output [SIZE - 1:0] out13,
    output [SIZE - 1:0] out14,
    output [SIZE - 1:0] out15,
    output [SIZE - 1:0] out16,
    output [SIZE - 1:0] out17,
    output [SIZE - 1:0] out18,
    output [SIZE - 1:0] out19,
    output [SIZE - 1:0] out20,
    output [SIZE - 1:0] out21,
    output [SIZE - 1:0] out22,
    output [SIZE - 1:0] out23,
    output [SIZE - 1:0] out24,
    output [SIZE - 1:0] out25,
    output [SIZE - 1:0] out26,
    output [SIZE - 1:0] out27,
    output [SIZE - 1:0] out28,
    output [SIZE - 1:0] out29,
    output [SIZE - 1:0] out30,
    output [SIZE - 1:0] out31,
    output [SIZE - 1:0] out32,
    output [SIZE - 1:0] out33,
    output [SIZE - 1:0] out34,
    output [SIZE - 1:0] out35,
    output [SIZE - 1:0] out36,
    output [SIZE - 1:0] out37,
    output [SIZE - 1:0] out38,
    output [SIZE - 1:0] out39,
    output [SIZE - 1:0] out40,
    output [SIZE - 1:0] out41,
    output [SIZE - 1:0] out42,
    output [SIZE - 1:0] out43,
    output [SIZE - 1:0] out44,
    output [SIZE - 1:0] out45,
    output [SIZE - 1:0] out46,
    output [SIZE - 1:0] out47,
    output [SIZE - 1:0] out48,
    output [SIZE - 1:0] out49,
    output [SIZE - 1:0] out50,
    output [SIZE - 1:0] out51,
    output [SIZE - 1:0] out52,
    output [SIZE - 1:0] out53,
    output [SIZE - 1:0] out54,
    output [SIZE - 1:0] out55,
    output [SIZE - 1:0] out56,
    output [SIZE - 1:0] out57,
    output [SIZE - 1:0] out58,
    output [SIZE - 1:0] out59,
    output [SIZE - 1:0] out60,
    output [SIZE - 1:0] out61,
    output [SIZE - 1:0] out62,
    output [SIZE - 1:0] out63,
    output [SIZE - 1:0] out64,
    output [SIZE - 1:0] out65,
    output [SIZE - 1:0] out66,
    output [SIZE - 1:0] out67,
    output [SIZE - 1:0] out68,
    output [SIZE - 1:0] out69,
    output [SIZE - 1:0] out70,
    output [SIZE - 1:0] out71,
    output [SIZE - 1:0] out72,
    output [SIZE - 1:0] out73,
    output [SIZE - 1:0] out74,
    output [SIZE - 1:0] out75,
    output [SIZE - 1:0] out76,
    output [SIZE - 1:0] out77,
    output [SIZE - 1:0] out78,
    output [SIZE - 1:0] out79,
    output [SIZE - 1:0] out80,
    output [SIZE - 1:0] out81,
    output [SIZE - 1:0] out82,
    output [SIZE - 1:0] out83,
    output [SIZE - 1:0] out84,
    output [SIZE - 1:0] out85,
    output [SIZE - 1:0] out86,
    output [SIZE - 1:0] out87,
    output [SIZE - 1:0] out88,
    output [SIZE - 1:0] out89,
    output [SIZE - 1:0] out90,
    output [SIZE - 1:0] out91,
    output [SIZE - 1:0] out92,
    output [SIZE - 1:0] out93,
    output [SIZE - 1:0] out94,
    output [SIZE - 1:0] out95,
    output [SIZE - 1:0] out96,
    output [SIZE - 1:0] out97,
    output [SIZE - 1:0] out98,
    output [SIZE - 1:0] out99,
    output [SIZE - 1:0] out100,
    output [SIZE - 1:0] out101,
    output [SIZE - 1:0] out102,
    output [SIZE - 1:0] out103,
    output [SIZE - 1:0] out104,
    output [SIZE - 1:0] out105,
    output [SIZE - 1:0] out106,
    output [SIZE - 1:0] out107,
    output [SIZE - 1:0] out108,
    output [SIZE - 1:0] out109,
    output [SIZE - 1:0] out110,
    output [SIZE - 1:0] out111,
    output [SIZE - 1:0] out112,
    output [SIZE - 1:0] out113,
    output [SIZE - 1:0] out114,
    output [SIZE - 1:0] out115,
    output [SIZE - 1:0] out116,
    output [SIZE - 1:0] out117,
    output [SIZE - 1:0] out118,
    output [SIZE - 1:0] out119,
    output [SIZE - 1:0] out120,
    output [SIZE - 1:0] out121,
    output [SIZE - 1:0] out122,
    output [SIZE - 1:0] out123,
    output [SIZE - 1:0] out124,
    output [SIZE - 1:0] out125,
    output [SIZE - 1:0] out126,
    output [SIZE - 1:0] out127,
    output [SIZE - 1:0] out128,
    output [SIZE - 1:0] out129,
    output [SIZE - 1:0] out130,
    output [SIZE - 1:0] out131,
    output [SIZE - 1:0] out132,
    output [SIZE - 1:0] out133,
    output [SIZE - 1:0] out134,
    output [SIZE - 1:0] out135,
    output [SIZE - 1:0] out136,
    output [SIZE - 1:0] out137,
    output [SIZE - 1:0] out138,
    output [SIZE - 1:0] out139,
    output [SIZE - 1:0] out140,
    output [SIZE - 1:0] out141,
    output [SIZE - 1:0] out142,
    output [SIZE - 1:0] out143,
    output [SIZE - 1:0] out144,
    output [SIZE - 1:0] out145,
    output [SIZE - 1:0] out146,
    output [SIZE - 1:0] out147,
    output [SIZE - 1:0] out148,
    output [SIZE - 1:0] out149,
    output [SIZE - 1:0] out150,
    output [SIZE - 1:0] out151,
    output [SIZE - 1:0] out152,
    output [SIZE - 1:0] out153,
    output [SIZE - 1:0] out154,
    output [SIZE - 1:0] out155,
    output [SIZE - 1:0] out156,
    output [SIZE - 1:0] out157,
    output [SIZE - 1:0] out158,
    output [SIZE - 1:0] out159,
    output [SIZE - 1:0] out160,
    output [SIZE - 1:0] out161,
    output [SIZE - 1:0] out162,
    output [SIZE - 1:0] out163,
    output [SIZE - 1:0] out164,
    output [SIZE - 1:0] out165,
    output [SIZE - 1:0] out166,
    output [SIZE - 1:0] out167,
    output [SIZE - 1:0] out168,
    output [SIZE - 1:0] out169,
    output [SIZE - 1:0] out170,
    output [SIZE - 1:0] out171,
    output [SIZE - 1:0] out172,
    output [SIZE - 1:0] out173,
    output [SIZE - 1:0] out174,
    output [SIZE - 1:0] out175,
    output [SIZE - 1:0] out176,
    output [SIZE - 1:0] out177,
    output [SIZE - 1:0] out178,
    output [SIZE - 1:0] out179,
    output [SIZE - 1:0] out180,
    output [SIZE - 1:0] out181,
    output [SIZE - 1:0] out182,
    output [SIZE - 1:0] out183,
    output [SIZE - 1:0] out184,
    output [SIZE - 1:0] out185,
    output [SIZE - 1:0] out186,
    output [SIZE - 1:0] out187,
    output [SIZE - 1:0] out188,
    output [SIZE - 1:0] out189,
    output [SIZE - 1:0] out190,
    output [SIZE - 1:0] out191,
    output [SIZE - 1:0] out192,
    output [SIZE - 1:0] out193,
    output [SIZE - 1:0] out194,
    output [SIZE - 1:0] out195,
    output [SIZE - 1:0] out196,
    output [SIZE - 1:0] out197,
    output [SIZE - 1:0] out198,
    output [SIZE - 1:0] out199,
    output [SIZE - 1:0] out200,
    output [SIZE - 1:0] out201,
    output [SIZE - 1:0] out202,
    output [SIZE - 1:0] out203,
    output [SIZE - 1:0] out204,
    output [SIZE - 1:0] out205,
    output [SIZE - 1:0] out206,
    output [SIZE - 1:0] out207,
    output [SIZE - 1:0] out208,
    output [SIZE - 1:0] out209,
    output [SIZE - 1:0] out210,
    output [SIZE - 1:0] out211,
    output [SIZE - 1:0] out212,
    output [SIZE - 1:0] out213,
    output [SIZE - 1:0] out214,
    output [SIZE - 1:0] out215,
    output [SIZE - 1:0] out216,
    output [SIZE - 1:0] out217,
    output [SIZE - 1:0] out218,
    output [SIZE - 1:0] out219,
    output [SIZE - 1:0] out220,
    output [SIZE - 1:0] out221,
    output [SIZE - 1:0] out222,
    output [SIZE - 1:0] out223,
    output [SIZE - 1:0] out224,
    output [SIZE - 1:0] out225,
    output [SIZE - 1:0] out226,
    output [SIZE - 1:0] out227,
    output [SIZE - 1:0] out228,
    output [SIZE - 1:0] out229,
    output [SIZE - 1:0] out230,
    output [SIZE - 1:0] out231,
    output [SIZE - 1:0] out232,
    output [SIZE - 1:0] out233,
    output [SIZE - 1:0] out234,
    output [SIZE - 1:0] out235,
    output [SIZE - 1:0] out236,
    output [SIZE - 1:0] out237,
    output [SIZE - 1:0] out238,
    output [SIZE - 1:0] out239,
    output [SIZE - 1:0] out240,
    output [SIZE - 1:0] out241,
    output [SIZE - 1:0] out242,
    output [SIZE - 1:0] out243,
    output [SIZE - 1:0] out244,
    output [SIZE - 1:0] out245,
    output [SIZE - 1:0] out246,
    output [SIZE - 1:0] out247,
    output [SIZE - 1:0] out248,
    output [SIZE - 1:0] out249,
    output [SIZE - 1:0] out250,
    output [SIZE - 1:0] out251,
    output [SIZE - 1:0] out252,
    output [SIZE - 1:0] out253,
    output [SIZE - 1:0] out254,
    output [SIZE - 1:0] out255,
    output [SIZE - 1:0] out256,
    output [SIZE - 1:0] out257,
    output [SIZE - 1:0] out258,
    output [SIZE - 1:0] out259,
    output [SIZE - 1:0] out260,
    output [SIZE - 1:0] out261,
    output [SIZE - 1:0] out262,
    output [SIZE - 1:0] out263,
    output [SIZE - 1:0] out264,
    output [SIZE - 1:0] out265,
    output [SIZE - 1:0] out266,
    output [SIZE - 1:0] out267,
    output [SIZE - 1:0] out268,
    output [SIZE - 1:0] out269,
    output [SIZE - 1:0] out270,
    output [SIZE - 1:0] out271,
    output [SIZE - 1:0] out272,
    output [SIZE - 1:0] out273,
    output [SIZE - 1:0] out274,
    output [SIZE - 1:0] out275,
    output [SIZE - 1:0] out276,
    output [SIZE - 1:0] out277,
    output [SIZE - 1:0] out278,
    output [SIZE - 1:0] out279,
    output [SIZE - 1:0] out280,
    output [SIZE - 1:0] out281,
    output [SIZE - 1:0] out282,
    output [SIZE - 1:0] out283,
    output [SIZE - 1:0] out284,
    output [SIZE - 1:0] out285,
    output [SIZE - 1:0] out286,
    output [SIZE - 1:0] out287,
    output [SIZE - 1:0] out288,
    output [SIZE - 1:0] out289,
    output [SIZE - 1:0] out290,
    output [SIZE - 1:0] out291,
    output [SIZE - 1:0] out292,
    output [SIZE - 1:0] out293,
    output [SIZE - 1:0] out294,
    output [SIZE - 1:0] out295,
    output [SIZE - 1:0] out296,
    output [SIZE - 1:0] out297,
    output [SIZE - 1:0] out298,
    output [SIZE - 1:0] out299,
    output [SIZE - 1:0] out300,
    output [SIZE - 1:0] out301,
    output [SIZE - 1:0] out302,
    output [SIZE - 1:0] out303,
    output [SIZE - 1:0] out304,
    output [SIZE - 1:0] out305,
    output [SIZE - 1:0] out306,
    output [SIZE - 1:0] out307,
    output [SIZE - 1:0] out308,
    output [SIZE - 1:0] out309,
    output [SIZE - 1:0] out310,
    output [SIZE - 1:0] out311,
    output [SIZE - 1:0] out312,
    output [SIZE - 1:0] out313,
    output [SIZE - 1:0] out314,
    output [SIZE - 1:0] out315,
    output [SIZE - 1:0] out316,
    output [SIZE - 1:0] out317,
    output [SIZE - 1:0] out318,
    output [SIZE - 1:0] out319,
    output [SIZE - 1:0] out320,
    output [SIZE - 1:0] out321,
    output [SIZE - 1:0] out322,
    output [SIZE - 1:0] out323,
    output [SIZE - 1:0] out324,
    output [SIZE - 1:0] out325,
    output [SIZE - 1:0] out326,
    output [SIZE - 1:0] out327,
    output [SIZE - 1:0] out328,
    output [SIZE - 1:0] out329,
    output [SIZE - 1:0] out330,
    output [SIZE - 1:0] out331,
    output [SIZE - 1:0] out332,
    output [SIZE - 1:0] out333,
    output [SIZE - 1:0] out334,
    output [SIZE - 1:0] out335,
    output [SIZE - 1:0] out336,
    output [SIZE - 1:0] out337,
    output [SIZE - 1:0] out338,
    output [SIZE - 1:0] out339,
    output [SIZE - 1:0] out340,
    output [SIZE - 1:0] out341,
    output [SIZE - 1:0] out342,
    output [SIZE - 1:0] out343,
    output [SIZE - 1:0] out344,
    output [SIZE - 1:0] out345,
    output [SIZE - 1:0] out346,
    output [SIZE - 1:0] out347,
    output [SIZE - 1:0] out348,
    output [SIZE - 1:0] out349,
    output [SIZE - 1:0] out350,
    output [SIZE - 1:0] out351,
    output [SIZE - 1:0] out352,
    output [SIZE - 1:0] out353,
    output [SIZE - 1:0] out354,
    output [SIZE - 1:0] out355,
    output [SIZE - 1:0] out356,
    output [SIZE - 1:0] out357,
    output [SIZE - 1:0] out358,
    output [SIZE - 1:0] out359,
    output [SIZE - 1:0] out360,
    output [SIZE - 1:0] out361,
    output [SIZE - 1:0] out362,
    output [SIZE - 1:0] out363,
    output [SIZE - 1:0] out364,
    output [SIZE - 1:0] out365,
    output [SIZE - 1:0] out366,
    output [SIZE - 1:0] out367,
    output [SIZE - 1:0] out368,
    output [SIZE - 1:0] out369,
    output [SIZE - 1:0] out370,
    output [SIZE - 1:0] out371,
    output [SIZE - 1:0] out372,
    output [SIZE - 1:0] out373,
    output [SIZE - 1:0] out374,
    output [SIZE - 1:0] out375,
    output [SIZE - 1:0] out376,
    output [SIZE - 1:0] out377,
    output [SIZE - 1:0] out378,
    output [SIZE - 1:0] out379,
    output [SIZE - 1:0] out380,
    output [SIZE - 1:0] out381,
    output [SIZE - 1:0] out382,
    output [SIZE - 1:0] out383,
    output [SIZE - 1:0] out384,
    output [SIZE - 1:0] out385,
    output [SIZE - 1:0] out386,
    output [SIZE - 1:0] out387,
    output [SIZE - 1:0] out388,
    output [SIZE - 1:0] out389,
    output [SIZE - 1:0] out390,
    output [SIZE - 1:0] out391,
    output [SIZE - 1:0] out392,
    output [SIZE - 1:0] out393,
    output [SIZE - 1:0] out394,
    output [SIZE - 1:0] out395,
    output [SIZE - 1:0] out396,
    output [SIZE - 1:0] out397,
    output [SIZE - 1:0] out398,
    output [SIZE - 1:0] out399,
    output [SIZE - 1:0] out400,
    output [SIZE - 1:0] out401,
    output [SIZE - 1:0] out402,
    output [SIZE - 1:0] out403,
    output [SIZE - 1:0] out404,
    output [SIZE - 1:0] out405,
    output [SIZE - 1:0] out406,
    output [SIZE - 1:0] out407,
    output [SIZE - 1:0] out408,
    output [SIZE - 1:0] out409,
    output [SIZE - 1:0] out410,
    output [SIZE - 1:0] out411,
    output [SIZE - 1:0] out412,
    output [SIZE - 1:0] out413,
    output [SIZE - 1:0] out414,
    output [SIZE - 1:0] out415,
    output [SIZE - 1:0] out416,
    output [SIZE - 1:0] out417,
    output [SIZE - 1:0] out418,
    output [SIZE - 1:0] out419,
    output [SIZE - 1:0] out420,
    output [SIZE - 1:0] out421,
    output [SIZE - 1:0] out422,
    output [SIZE - 1:0] out423,
    output [SIZE - 1:0] out424,
    output [SIZE - 1:0] out425,
    output [SIZE - 1:0] out426,
    output [SIZE - 1:0] out427,
    output [SIZE - 1:0] out428,
    output [SIZE - 1:0] out429,
    output [SIZE - 1:0] out430,
    output [SIZE - 1:0] out431,
    output [SIZE - 1:0] out432,
    output [SIZE - 1:0] out433,
    output [SIZE - 1:0] out434,
    output [SIZE - 1:0] out435,
    output [SIZE - 1:0] out436,
    output [SIZE - 1:0] out437,
    output [SIZE - 1:0] out438,
    output [SIZE - 1:0] out439,
    output [SIZE - 1:0] out440,
    output [SIZE - 1:0] out441,
    output [SIZE - 1:0] out442,
    output [SIZE - 1:0] out443,
    output [SIZE - 1:0] out444,
    output [SIZE - 1:0] out445,
    output [SIZE - 1:0] out446,
    output [SIZE - 1:0] out447,
    output [SIZE - 1:0] out448,
    output [SIZE - 1:0] out449,
    output [SIZE - 1:0] out450,
    output [SIZE - 1:0] out451,
    output [SIZE - 1:0] out452,
    output [SIZE - 1:0] out453,
    output [SIZE - 1:0] out454,
    output [SIZE - 1:0] out455,
    output [SIZE - 1:0] out456,
    output [SIZE - 1:0] out457,
    output [SIZE - 1:0] out458,
    output [SIZE - 1:0] out459,
    output [SIZE - 1:0] out460,
    output [SIZE - 1:0] out461,
    output [SIZE - 1:0] out462,
    output [SIZE - 1:0] out463,
    output [SIZE - 1:0] out464,
    output [SIZE - 1:0] out465,
    output [SIZE - 1:0] out466,
    output [SIZE - 1:0] out467,
    output [SIZE - 1:0] out468,
    output [SIZE - 1:0] out469,
    output [SIZE - 1:0] out470,
    output [SIZE - 1:0] out471,
    output [SIZE - 1:0] out472,
    output [SIZE - 1:0] out473,
    output [SIZE - 1:0] out474,
    output [SIZE - 1:0] out475,
    output [SIZE - 1:0] out476,
    output [SIZE - 1:0] out477,
    output [SIZE - 1:0] out478,
    output [SIZE - 1:0] out479,
    output [SIZE - 1:0] out480,
    output [SIZE - 1:0] out481,
    output [SIZE - 1:0] out482,
    output [SIZE - 1:0] out483,
    output [SIZE - 1:0] out484,
    output [SIZE - 1:0] out485,
    output [SIZE - 1:0] out486,
    output [SIZE - 1:0] out487,
    output [SIZE - 1:0] out488,
    output [SIZE - 1:0] out489,
    output [SIZE - 1:0] out490,
    output [SIZE - 1:0] out491,
    output [SIZE - 1:0] out492,
    output [SIZE - 1:0] out493,
    output [SIZE - 1:0] out494,
    output [SIZE - 1:0] out495,
    output [SIZE - 1:0] out496,
    output [SIZE - 1:0] out497,
    output [SIZE - 1:0] out498,
    output [SIZE - 1:0] out499,
    output [SIZE - 1:0] out500,
    output [SIZE - 1:0] out501,
    output [SIZE - 1:0] out502,
    output [SIZE - 1:0] out503,
    output [SIZE - 1:0] out504,
    output [SIZE - 1:0] out505,
    output [SIZE - 1:0] out506,
    output [SIZE - 1:0] out507,
    output [SIZE - 1:0] out508,
    output [SIZE - 1:0] out509,
    output [SIZE - 1:0] out510,
    output [SIZE - 1:0] out511,
    output [SIZE - 1:0] out512,
    output [SIZE - 1:0] out513,
    output [SIZE - 1:0] out514,
    output [SIZE - 1:0] out515,
    output [SIZE - 1:0] out516,
    output [SIZE - 1:0] out517,
    output [SIZE - 1:0] out518,
    output [SIZE - 1:0] out519,
    output [SIZE - 1:0] out520,
    output [SIZE - 1:0] out521,
    output [SIZE - 1:0] out522,
    output [SIZE - 1:0] out523,
    output [SIZE - 1:0] out524,
    output [SIZE - 1:0] out525,
    output [SIZE - 1:0] out526,
    output [SIZE - 1:0] out527,
    output [SIZE - 1:0] out528,
    output [SIZE - 1:0] out529,
    output [SIZE - 1:0] out530,
    output [SIZE - 1:0] out531,
    output [SIZE - 1:0] out532,
    output [SIZE - 1:0] out533,
    output [SIZE - 1:0] out534,
    output [SIZE - 1:0] out535,
    output [SIZE - 1:0] out536,
    output [SIZE - 1:0] out537,
    output [SIZE - 1:0] out538,
    output [SIZE - 1:0] out539,
    output [SIZE - 1:0] out540,
    output [SIZE - 1:0] out541,
    output [SIZE - 1:0] out542,
    output [SIZE - 1:0] out543,
    output [SIZE - 1:0] out544,
    output [SIZE - 1:0] out545,
    output [SIZE - 1:0] out546,
    output [SIZE - 1:0] out547,
    output [SIZE - 1:0] out548,
    output [SIZE - 1:0] out549,
    output [SIZE - 1:0] out550,
    output [SIZE - 1:0] out551,
    output [SIZE - 1:0] out552,
    output [SIZE - 1:0] out553,
    output [SIZE - 1:0] out554,
    output [SIZE - 1:0] out555,
    output [SIZE - 1:0] out556,
    output [SIZE - 1:0] out557,
    output [SIZE - 1:0] out558,
    output [SIZE - 1:0] out559,
    output [SIZE - 1:0] out560,
    output [SIZE - 1:0] out561,
    output [SIZE - 1:0] out562,
    output [SIZE - 1:0] out563,
    output [SIZE - 1:0] out564,
    output [SIZE - 1:0] out565,
    output [SIZE - 1:0] out566,
    output [SIZE - 1:0] out567,
    output [SIZE - 1:0] out568,
    output [SIZE - 1:0] out569,
    output [SIZE - 1:0] out570,
    output [SIZE - 1:0] out571,
    output [SIZE - 1:0] out572,
    output [SIZE - 1:0] out573,
    output [SIZE - 1:0] out574,
    output [SIZE - 1:0] out575,
    output [SIZE - 1:0] out576,
    output [SIZE - 1:0] out577,
    output [SIZE - 1:0] out578,
    output [SIZE - 1:0] out579,
    output [SIZE - 1:0] out580,
    output [SIZE - 1:0] out581,
    output [SIZE - 1:0] out582,
    output [SIZE - 1:0] out583,
    output [SIZE - 1:0] out584,
    output [SIZE - 1:0] out585,
    output [SIZE - 1:0] out586,
    output [SIZE - 1:0] out587,
    output [SIZE - 1:0] out588,
    output [SIZE - 1:0] out589,
    output [SIZE - 1:0] out590,
    output [SIZE - 1:0] out591,
    output [SIZE - 1:0] out592,
    output [SIZE - 1:0] out593,
    output [SIZE - 1:0] out594,
    output [SIZE - 1:0] out595,
    output [SIZE - 1:0] out596,
    output [SIZE - 1:0] out597,
    output [SIZE - 1:0] out598,
    output [SIZE - 1:0] out599,
    output [SIZE - 1:0] out600,
    output [SIZE - 1:0] out601,
    output [SIZE - 1:0] out602,
    output [SIZE - 1:0] out603,
    output [SIZE - 1:0] out604,
    output [SIZE - 1:0] out605,
    output [SIZE - 1:0] out606,
    output [SIZE - 1:0] out607,
    output [SIZE - 1:0] out608,
    output [SIZE - 1:0] out609,
    output [SIZE - 1:0] out610,
    output [SIZE - 1:0] out611,
    output [SIZE - 1:0] out612,
    output [SIZE - 1:0] out613,
    output [SIZE - 1:0] out614,
    output [SIZE - 1:0] out615,
    output [SIZE - 1:0] out616,
    output [SIZE - 1:0] out617,
    output [SIZE - 1:0] out618,
    output [SIZE - 1:0] out619,
    output [SIZE - 1:0] out620,
    output [SIZE - 1:0] out621,
    output [SIZE - 1:0] out622,
    output [SIZE - 1:0] out623,
    output [SIZE - 1:0] out624,
    output [SIZE - 1:0] out625,
    output [SIZE - 1:0] out626,
    output [SIZE - 1:0] out627,
    output [SIZE - 1:0] out628,
    output [SIZE - 1:0] out629,
    output [SIZE - 1:0] out630,
    output [SIZE - 1:0] out631,
    output [SIZE - 1:0] out632,
    output [SIZE - 1:0] out633,
    output [SIZE - 1:0] out634,
    output [SIZE - 1:0] out635,
    output [SIZE - 1:0] out636,
    output [SIZE - 1:0] out637,
    output [SIZE - 1:0] out638,
    output [SIZE - 1:0] out639,
    output [SIZE - 1:0] out640,
    output [SIZE - 1:0] out641,
    output [SIZE - 1:0] out642,
    output [SIZE - 1:0] out643,
    output [SIZE - 1:0] out644,
    output [SIZE - 1:0] out645,
    output [SIZE - 1:0] out646,
    output [SIZE - 1:0] out647,
    output [SIZE - 1:0] out648,
    output [SIZE - 1:0] out649,
    output [SIZE - 1:0] out650,
    output [SIZE - 1:0] out651,
    output [SIZE - 1:0] out652,
    output [SIZE - 1:0] out653,
    output [SIZE - 1:0] out654,
    output [SIZE - 1:0] out655,
    output [SIZE - 1:0] out656,
    output [SIZE - 1:0] out657,
    output [SIZE - 1:0] out658,
    output [SIZE - 1:0] out659,
    output [SIZE - 1:0] out660,
    output [SIZE - 1:0] out661,
    output [SIZE - 1:0] out662,
    output [SIZE - 1:0] out663,
    output [SIZE - 1:0] out664,
    output [SIZE - 1:0] out665,
    output [SIZE - 1:0] out666,
    output [SIZE - 1:0] out667,
    output [SIZE - 1:0] out668,
    output [SIZE - 1:0] out669,
    output [SIZE - 1:0] out670,
    output [SIZE - 1:0] out671,
    output [SIZE - 1:0] out672,
    output [SIZE - 1:0] out673,
    output [SIZE - 1:0] out674,
    output [SIZE - 1:0] out675,
    output [SIZE - 1:0] out676,
    output [SIZE - 1:0] out677,
    output [SIZE - 1:0] out678,
    output [SIZE - 1:0] out679,
    output [SIZE - 1:0] out680,
    output [SIZE - 1:0] out681,
    output [SIZE - 1:0] out682,
    output [SIZE - 1:0] out683,
    output [SIZE - 1:0] out684,
    output [SIZE - 1:0] out685,
    output [SIZE - 1:0] out686,
    output [SIZE - 1:0] out687,
    output [SIZE - 1:0] out688,
    output [SIZE - 1:0] out689,
    output [SIZE - 1:0] out690,
    output [SIZE - 1:0] out691,
    output [SIZE - 1:0] out692,
    output [SIZE - 1:0] out693,
    output [SIZE - 1:0] out694,
    output [SIZE - 1:0] out695,
    output [SIZE - 1:0] out696,
    output [SIZE - 1:0] out697,
    output [SIZE - 1:0] out698,
    output [SIZE - 1:0] out699,
    output [SIZE - 1:0] out700,
    output [SIZE - 1:0] out701,
    output [SIZE - 1:0] out702,
    output [SIZE - 1:0] out703,
    output [SIZE - 1:0] out704,
    output [SIZE - 1:0] out705,
    output [SIZE - 1:0] out706,
    output [SIZE - 1:0] out707,
    output [SIZE - 1:0] out708,
    output [SIZE - 1:0] out709,
    output [SIZE - 1:0] out710,
    output [SIZE - 1:0] out711,
    output [SIZE - 1:0] out712,
    output [SIZE - 1:0] out713,
    output [SIZE - 1:0] out714,
    output [SIZE - 1:0] out715,
    output [SIZE - 1:0] out716,
    output [SIZE - 1:0] out717,
    output [SIZE - 1:0] out718,
    output [SIZE - 1:0] out719,
    output [SIZE - 1:0] out720,
    output [SIZE - 1:0] out721,
    output [SIZE - 1:0] out722,
    output [SIZE - 1:0] out723,
    output [SIZE - 1:0] out724,
    output [SIZE - 1:0] out725,
    output [SIZE - 1:0] out726,
    output [SIZE - 1:0] out727,
    output [SIZE - 1:0] out728,
    output [SIZE - 1:0] out729,
    output [SIZE - 1:0] out730,
    output [SIZE - 1:0] out731,
    output [SIZE - 1:0] out732,
    output [SIZE - 1:0] out733,
    output [SIZE - 1:0] out734,
    output [SIZE - 1:0] out735,
    output [SIZE - 1:0] out736,
    output [SIZE - 1:0] out737,
    output [SIZE - 1:0] out738,
    output [SIZE - 1:0] out739,
    output [SIZE - 1:0] out740,
    output [SIZE - 1:0] out741,
    output [SIZE - 1:0] out742,
    output [SIZE - 1:0] out743,
    output [SIZE - 1:0] out744,
    output [SIZE - 1:0] out745,
    output [SIZE - 1:0] out746,
    output [SIZE - 1:0] out747,
    output [SIZE - 1:0] out748,
    output [SIZE - 1:0] out749,
    output [SIZE - 1:0] out750,
    output [SIZE - 1:0] out751,
    output [SIZE - 1:0] out752,
    output [SIZE - 1:0] out753,
    output [SIZE - 1:0] out754,
    output [SIZE - 1:0] out755,
    output [SIZE - 1:0] out756,
    output [SIZE - 1:0] out757,
    output [SIZE - 1:0] out758,
    output [SIZE - 1:0] out759,
    output [SIZE - 1:0] out760,
    output [SIZE - 1:0] out761,
    output [SIZE - 1:0] out762,
    output [SIZE - 1:0] out763,
    output [SIZE - 1:0] out764,
    output [SIZE - 1:0] out765,
    output [SIZE - 1:0] out766,
    output [SIZE - 1:0] out767,
    output [SIZE - 1:0] out768,
    output [SIZE - 1:0] out769,
    output [SIZE - 1:0] out770,
    output [SIZE - 1:0] out771,
    output [SIZE - 1:0] out772,
    output [SIZE - 1:0] out773,
    output [SIZE - 1:0] out774,
    output [SIZE - 1:0] out775,
    output [SIZE - 1:0] out776,
    output [SIZE - 1:0] out777,
    output [SIZE - 1:0] out778,
    output [SIZE - 1:0] out779,
    output [SIZE - 1:0] out780,
    output [SIZE - 1:0] out781,
    output [SIZE - 1:0] out782,
    output [SIZE - 1:0] out783,
    output [SIZE - 1:0] out784,
    output [SIZE - 1:0] out785,
    output [SIZE - 1:0] out786,
    output [SIZE - 1:0] out787,
    output [SIZE - 1:0] out788,
    output [SIZE - 1:0] out789,
    output [SIZE - 1:0] out790,
    output [SIZE - 1:0] out791,
    output [SIZE - 1:0] out792,
    output [SIZE - 1:0] out793,
    output [SIZE - 1:0] out794,
    output [SIZE - 1:0] out795,
    output [SIZE - 1:0] out796,
    output [SIZE - 1:0] out797,
    output [SIZE - 1:0] out798,
    output [SIZE - 1:0] out799,
    output [SIZE - 1:0] out800,
    output [SIZE - 1:0] out801,
    output [SIZE - 1:0] out802,
    output [SIZE - 1:0] out803,
    output [SIZE - 1:0] out804,
    output [SIZE - 1:0] out805,
    output [SIZE - 1:0] out806,
    output [SIZE - 1:0] out807,
    output [SIZE - 1:0] out808,
    output [SIZE - 1:0] out809,
    output [SIZE - 1:0] out810,
    output [SIZE - 1:0] out811,
    output [SIZE - 1:0] out812,
    output [SIZE - 1:0] out813,
    output [SIZE - 1:0] out814,
    output [SIZE - 1:0] out815,
    output [SIZE - 1:0] out816,
    output [SIZE - 1:0] out817,
    output [SIZE - 1:0] out818,
    output [SIZE - 1:0] out819,
    output [SIZE - 1:0] out820,
    output [SIZE - 1:0] out821,
    output [SIZE - 1:0] out822,
    output [SIZE - 1:0] out823,
    output [SIZE - 1:0] out824,
    output [SIZE - 1:0] out825,
    output [SIZE - 1:0] out826,
    output [SIZE - 1:0] out827,
    output [SIZE - 1:0] out828,
    output [SIZE - 1:0] out829,
    output [SIZE - 1:0] out830,
    output [SIZE - 1:0] out831,
    output [SIZE - 1:0] out832,
    output [SIZE - 1:0] out833,
    output [SIZE - 1:0] out834,
    output [SIZE - 1:0] out835,
    output [SIZE - 1:0] out836,
    output [SIZE - 1:0] out837,
    output [SIZE - 1:0] out838,
    output [SIZE - 1:0] out839,
    output [SIZE - 1:0] out840,
    output [SIZE - 1:0] out841,
    output [SIZE - 1:0] out842,
    output [SIZE - 1:0] out843,
    output [SIZE - 1:0] out844,
    output [SIZE - 1:0] out845,
    output [SIZE - 1:0] out846,
    output [SIZE - 1:0] out847,
    output [SIZE - 1:0] out848,
    output [SIZE - 1:0] out849,
    output [SIZE - 1:0] out850,
    output [SIZE - 1:0] out851,
    output [SIZE - 1:0] out852,
    output [SIZE - 1:0] out853,
    output [SIZE - 1:0] out854,
    output [SIZE - 1:0] out855,
    output [SIZE - 1:0] out856,
    output [SIZE - 1:0] out857,
    output [SIZE - 1:0] out858,
    output [SIZE - 1:0] out859,
    output [SIZE - 1:0] out860,
    output [SIZE - 1:0] out861,
    output [SIZE - 1:0] out862,
    output [SIZE - 1:0] out863,
    output [SIZE - 1:0] out864,
    output [SIZE - 1:0] out865,
    output [SIZE - 1:0] out866,
    output [SIZE - 1:0] out867,
    output [SIZE - 1:0] out868,
    output [SIZE - 1:0] out869,
    output [SIZE - 1:0] out870,
    output [SIZE - 1:0] out871,
    output [SIZE - 1:0] out872,
    output [SIZE - 1:0] out873,
    output [SIZE - 1:0] out874,
    output [SIZE - 1:0] out875,
    output [SIZE - 1:0] out876,
    output [SIZE - 1:0] out877,
    output [SIZE - 1:0] out878,
    output [SIZE - 1:0] out879,
    output [SIZE - 1:0] out880,
    output [SIZE - 1:0] out881,
    output [SIZE - 1:0] out882,
    output [SIZE - 1:0] out883,
    output [SIZE - 1:0] out884,
    output [SIZE - 1:0] out885,
    output [SIZE - 1:0] out886,
    output [SIZE - 1:0] out887,
    output [SIZE - 1:0] out888,
    output [SIZE - 1:0] out889,
    output [SIZE - 1:0] out890,
    output [SIZE - 1:0] out891,
    output [SIZE - 1:0] out892,
    output [SIZE - 1:0] out893,
    output [SIZE - 1:0] out894,
    output [SIZE - 1:0] out895,
    output [SIZE - 1:0] out896,
    output [SIZE - 1:0] out897,
    output [SIZE - 1:0] out898,
    output [SIZE - 1:0] out899,
    output [SIZE - 1:0] out900,
    output [SIZE - 1:0] out901,
    output [SIZE - 1:0] out902,
    output [SIZE - 1:0] out903,
    output [SIZE - 1:0] out904,
    output [SIZE - 1:0] out905,
    output [SIZE - 1:0] out906,
    output [SIZE - 1:0] out907,
    output [SIZE - 1:0] out908,
    output [SIZE - 1:0] out909,
    output [SIZE - 1:0] out910,
    output [SIZE - 1:0] out911,
    output [SIZE - 1:0] out912,
    output [SIZE - 1:0] out913,
    output [SIZE - 1:0] out914,
    output [SIZE - 1:0] out915,
    output [SIZE - 1:0] out916,
    output [SIZE - 1:0] out917,
    output [SIZE - 1:0] out918,
    output [SIZE - 1:0] out919,
    output [SIZE - 1:0] out920,
    output [SIZE - 1:0] out921,
    output [SIZE - 1:0] out922,
    output [SIZE - 1:0] out923,
    output [SIZE - 1:0] out924,
    output [SIZE - 1:0] out925,
    output [SIZE - 1:0] out926,
    output [SIZE - 1:0] out927,
    output [SIZE - 1:0] out928,
    output [SIZE - 1:0] out929,
    output [SIZE - 1:0] out930,
    output [SIZE - 1:0] out931,
    output [SIZE - 1:0] out932,
    output [SIZE - 1:0] out933,
    output [SIZE - 1:0] out934,
    output [SIZE - 1:0] out935,
    output [SIZE - 1:0] out936,
    output [SIZE - 1:0] out937,
    output [SIZE - 1:0] out938,
    output [SIZE - 1:0] out939,
    output [SIZE - 1:0] out940,
    output [SIZE - 1:0] out941,
    output [SIZE - 1:0] out942,
    output [SIZE - 1:0] out943,
    output [SIZE - 1:0] out944,
    output [SIZE - 1:0] out945,
    output [SIZE - 1:0] out946,
    output [SIZE - 1:0] out947,
    output [SIZE - 1:0] out948,
    output [SIZE - 1:0] out949,
    output [SIZE - 1:0] out950,
    output [SIZE - 1:0] out951,
    output [SIZE - 1:0] out952,
    output [SIZE - 1:0] out953,
    output [SIZE - 1:0] out954,
    output [SIZE - 1:0] out955,
    output [SIZE - 1:0] out956,
    output [SIZE - 1:0] out957,
    output [SIZE - 1:0] out958,
    output [SIZE - 1:0] out959,
    output [SIZE - 1:0] out960,
    output [SIZE - 1:0] out961,
    output [SIZE - 1:0] out962,
    output [SIZE - 1:0] out963,
    output [SIZE - 1:0] out964,
    output [SIZE - 1:0] out965,
    output [SIZE - 1:0] out966,
    output [SIZE - 1:0] out967,
    output [SIZE - 1:0] out968,
    output [SIZE - 1:0] out969,
    output [SIZE - 1:0] out970,
    output [SIZE - 1:0] out971,
    output [SIZE - 1:0] out972,
    output [SIZE - 1:0] out973,
    output [SIZE - 1:0] out974,
    output [SIZE - 1:0] out975,
    output [SIZE - 1:0] out976,
    output [SIZE - 1:0] out977,
    output [SIZE - 1:0] out978,
    output [SIZE - 1:0] out979,
    output [SIZE - 1:0] out980,
    output [SIZE - 1:0] out981,
    output [SIZE - 1:0] out982,
    output [SIZE - 1:0] out983,
    output [SIZE - 1:0] out984,
    output [SIZE - 1:0] out985,
    output [SIZE - 1:0] out986,
    output [SIZE - 1:0] out987,
    output [SIZE - 1:0] out988,
    output [SIZE - 1:0] out989,
    output [SIZE - 1:0] out990,
    output [SIZE - 1:0] out991,
    output [SIZE - 1:0] out992,
    output [SIZE - 1:0] out993,
    output [SIZE - 1:0] out994,
    output [SIZE - 1:0] out995,
    output [SIZE - 1:0] out996,
    output [SIZE - 1:0] out997,
    output [SIZE - 1:0] out998,
    output [SIZE - 1:0] out999,
    output [SIZE - 1:0] out1000,
    output [SIZE - 1:0] out1001,
    output [SIZE - 1:0] out1002,
    output [SIZE - 1:0] out1003,
    output [SIZE - 1:0] out1004,
    output [SIZE - 1:0] out1005,
    output [SIZE - 1:0] out1006,
    output [SIZE - 1:0] out1007,
    output [SIZE - 1:0] out1008,
    output [SIZE - 1:0] out1009,
    output [SIZE - 1:0] out1010,
    output [SIZE - 1:0] out1011,
    output [SIZE - 1:0] out1012,
    output [SIZE - 1:0] out1013,
    output [SIZE - 1:0] out1014,
    output [SIZE - 1:0] out1015,
    output [SIZE - 1:0] out1016,
    output [SIZE - 1:0] out1017,
    output [SIZE - 1:0] out1018,
    output [SIZE - 1:0] out1019,
    output [SIZE - 1:0] out1020,
    output [SIZE - 1:0] out1021,
    output [SIZE - 1:0] out1022,
    output [SIZE - 1:0] out1023
);
    integer x, y, z;
    genvar i,j;

    reg [SIZE - 1:0] tmp [N - 1:0][STEP:0][1:0];
    wire [SIZE - 1:0] w [N - 1:0][STEP - 1:0][1:0];
    reg [3:0] stage;
    reg [3:0] counter;
    reg done;

    always@(*)begin
        tmp[0][0][0] = in0;
        tmp[1][0][0] = in1;
        tmp[2][0][0] = in2;
        tmp[3][0][0] = in3;
        tmp[4][0][0] = in4;
        tmp[5][0][0] = in5;
        tmp[6][0][0] = in6;
        tmp[7][0][0] = in7;
        tmp[8][0][0] = in8;
        tmp[9][0][0] = in9;
        tmp[10][0][0] = in10;
        tmp[11][0][0] = in11;
        tmp[12][0][0] = in12;
        tmp[13][0][0] = in13;
        tmp[14][0][0] = in14;
        tmp[15][0][0] = in15;
        tmp[16][0][0] = in16;
        tmp[17][0][0] = in17;
        tmp[18][0][0] = in18;
        tmp[19][0][0] = in19;
        tmp[20][0][0] = in20;
        tmp[21][0][0] = in21;
        tmp[22][0][0] = in22;
        tmp[23][0][0] = in23;
        tmp[24][0][0] = in24;
        tmp[25][0][0] = in25;
        tmp[26][0][0] = in26;
        tmp[27][0][0] = in27;
        tmp[28][0][0] = in28;
        tmp[29][0][0] = in29;
        tmp[30][0][0] = in30;
        tmp[31][0][0] = in31;
        tmp[32][0][0] = in32;
        tmp[33][0][0] = in33;
        tmp[34][0][0] = in34;
        tmp[35][0][0] = in35;
        tmp[36][0][0] = in36;
        tmp[37][0][0] = in37;
        tmp[38][0][0] = in38;
        tmp[39][0][0] = in39;
        tmp[40][0][0] = in40;
        tmp[41][0][0] = in41;
        tmp[42][0][0] = in42;
        tmp[43][0][0] = in43;
        tmp[44][0][0] = in44;
        tmp[45][0][0] = in45;
        tmp[46][0][0] = in46;
        tmp[47][0][0] = in47;
        tmp[48][0][0] = in48;
        tmp[49][0][0] = in49;
        tmp[50][0][0] = in50;
        tmp[51][0][0] = in51;
        tmp[52][0][0] = in52;
        tmp[53][0][0] = in53;
        tmp[54][0][0] = in54;
        tmp[55][0][0] = in55;
        tmp[56][0][0] = in56;
        tmp[57][0][0] = in57;
        tmp[58][0][0] = in58;
        tmp[59][0][0] = in59;
        tmp[60][0][0] = in60;
        tmp[61][0][0] = in61;
        tmp[62][0][0] = in62;
        tmp[63][0][0] = in63;
        tmp[64][0][0] = in64;
        tmp[65][0][0] = in65;
        tmp[66][0][0] = in66;
        tmp[67][0][0] = in67;
        tmp[68][0][0] = in68;
        tmp[69][0][0] = in69;
        tmp[70][0][0] = in70;
        tmp[71][0][0] = in71;
        tmp[72][0][0] = in72;
        tmp[73][0][0] = in73;
        tmp[74][0][0] = in74;
        tmp[75][0][0] = in75;
        tmp[76][0][0] = in76;
        tmp[77][0][0] = in77;
        tmp[78][0][0] = in78;
        tmp[79][0][0] = in79;
        tmp[80][0][0] = in80;
        tmp[81][0][0] = in81;
        tmp[82][0][0] = in82;
        tmp[83][0][0] = in83;
        tmp[84][0][0] = in84;
        tmp[85][0][0] = in85;
        tmp[86][0][0] = in86;
        tmp[87][0][0] = in87;
        tmp[88][0][0] = in88;
        tmp[89][0][0] = in89;
        tmp[90][0][0] = in90;
        tmp[91][0][0] = in91;
        tmp[92][0][0] = in92;
        tmp[93][0][0] = in93;
        tmp[94][0][0] = in94;
        tmp[95][0][0] = in95;
        tmp[96][0][0] = in96;
        tmp[97][0][0] = in97;
        tmp[98][0][0] = in98;
        tmp[99][0][0] = in99;
        tmp[100][0][0] = in100;
        tmp[101][0][0] = in101;
        tmp[102][0][0] = in102;
        tmp[103][0][0] = in103;
        tmp[104][0][0] = in104;
        tmp[105][0][0] = in105;
        tmp[106][0][0] = in106;
        tmp[107][0][0] = in107;
        tmp[108][0][0] = in108;
        tmp[109][0][0] = in109;
        tmp[110][0][0] = in110;
        tmp[111][0][0] = in111;
        tmp[112][0][0] = in112;
        tmp[113][0][0] = in113;
        tmp[114][0][0] = in114;
        tmp[115][0][0] = in115;
        tmp[116][0][0] = in116;
        tmp[117][0][0] = in117;
        tmp[118][0][0] = in118;
        tmp[119][0][0] = in119;
        tmp[120][0][0] = in120;
        tmp[121][0][0] = in121;
        tmp[122][0][0] = in122;
        tmp[123][0][0] = in123;
        tmp[124][0][0] = in124;
        tmp[125][0][0] = in125;
        tmp[126][0][0] = in126;
        tmp[127][0][0] = in127;
        tmp[128][0][0] = in128;
        tmp[129][0][0] = in129;
        tmp[130][0][0] = in130;
        tmp[131][0][0] = in131;
        tmp[132][0][0] = in132;
        tmp[133][0][0] = in133;
        tmp[134][0][0] = in134;
        tmp[135][0][0] = in135;
        tmp[136][0][0] = in136;
        tmp[137][0][0] = in137;
        tmp[138][0][0] = in138;
        tmp[139][0][0] = in139;
        tmp[140][0][0] = in140;
        tmp[141][0][0] = in141;
        tmp[142][0][0] = in142;
        tmp[143][0][0] = in143;
        tmp[144][0][0] = in144;
        tmp[145][0][0] = in145;
        tmp[146][0][0] = in146;
        tmp[147][0][0] = in147;
        tmp[148][0][0] = in148;
        tmp[149][0][0] = in149;
        tmp[150][0][0] = in150;
        tmp[151][0][0] = in151;
        tmp[152][0][0] = in152;
        tmp[153][0][0] = in153;
        tmp[154][0][0] = in154;
        tmp[155][0][0] = in155;
        tmp[156][0][0] = in156;
        tmp[157][0][0] = in157;
        tmp[158][0][0] = in158;
        tmp[159][0][0] = in159;
        tmp[160][0][0] = in160;
        tmp[161][0][0] = in161;
        tmp[162][0][0] = in162;
        tmp[163][0][0] = in163;
        tmp[164][0][0] = in164;
        tmp[165][0][0] = in165;
        tmp[166][0][0] = in166;
        tmp[167][0][0] = in167;
        tmp[168][0][0] = in168;
        tmp[169][0][0] = in169;
        tmp[170][0][0] = in170;
        tmp[171][0][0] = in171;
        tmp[172][0][0] = in172;
        tmp[173][0][0] = in173;
        tmp[174][0][0] = in174;
        tmp[175][0][0] = in175;
        tmp[176][0][0] = in176;
        tmp[177][0][0] = in177;
        tmp[178][0][0] = in178;
        tmp[179][0][0] = in179;
        tmp[180][0][0] = in180;
        tmp[181][0][0] = in181;
        tmp[182][0][0] = in182;
        tmp[183][0][0] = in183;
        tmp[184][0][0] = in184;
        tmp[185][0][0] = in185;
        tmp[186][0][0] = in186;
        tmp[187][0][0] = in187;
        tmp[188][0][0] = in188;
        tmp[189][0][0] = in189;
        tmp[190][0][0] = in190;
        tmp[191][0][0] = in191;
        tmp[192][0][0] = in192;
        tmp[193][0][0] = in193;
        tmp[194][0][0] = in194;
        tmp[195][0][0] = in195;
        tmp[196][0][0] = in196;
        tmp[197][0][0] = in197;
        tmp[198][0][0] = in198;
        tmp[199][0][0] = in199;
        tmp[200][0][0] = in200;
        tmp[201][0][0] = in201;
        tmp[202][0][0] = in202;
        tmp[203][0][0] = in203;
        tmp[204][0][0] = in204;
        tmp[205][0][0] = in205;
        tmp[206][0][0] = in206;
        tmp[207][0][0] = in207;
        tmp[208][0][0] = in208;
        tmp[209][0][0] = in209;
        tmp[210][0][0] = in210;
        tmp[211][0][0] = in211;
        tmp[212][0][0] = in212;
        tmp[213][0][0] = in213;
        tmp[214][0][0] = in214;
        tmp[215][0][0] = in215;
        tmp[216][0][0] = in216;
        tmp[217][0][0] = in217;
        tmp[218][0][0] = in218;
        tmp[219][0][0] = in219;
        tmp[220][0][0] = in220;
        tmp[221][0][0] = in221;
        tmp[222][0][0] = in222;
        tmp[223][0][0] = in223;
        tmp[224][0][0] = in224;
        tmp[225][0][0] = in225;
        tmp[226][0][0] = in226;
        tmp[227][0][0] = in227;
        tmp[228][0][0] = in228;
        tmp[229][0][0] = in229;
        tmp[230][0][0] = in230;
        tmp[231][0][0] = in231;
        tmp[232][0][0] = in232;
        tmp[233][0][0] = in233;
        tmp[234][0][0] = in234;
        tmp[235][0][0] = in235;
        tmp[236][0][0] = in236;
        tmp[237][0][0] = in237;
        tmp[238][0][0] = in238;
        tmp[239][0][0] = in239;
        tmp[240][0][0] = in240;
        tmp[241][0][0] = in241;
        tmp[242][0][0] = in242;
        tmp[243][0][0] = in243;
        tmp[244][0][0] = in244;
        tmp[245][0][0] = in245;
        tmp[246][0][0] = in246;
        tmp[247][0][0] = in247;
        tmp[248][0][0] = in248;
        tmp[249][0][0] = in249;
        tmp[250][0][0] = in250;
        tmp[251][0][0] = in251;
        tmp[252][0][0] = in252;
        tmp[253][0][0] = in253;
        tmp[254][0][0] = in254;
        tmp[255][0][0] = in255;
        tmp[256][0][0] = in256;
        tmp[257][0][0] = in257;
        tmp[258][0][0] = in258;
        tmp[259][0][0] = in259;
        tmp[260][0][0] = in260;
        tmp[261][0][0] = in261;
        tmp[262][0][0] = in262;
        tmp[263][0][0] = in263;
        tmp[264][0][0] = in264;
        tmp[265][0][0] = in265;
        tmp[266][0][0] = in266;
        tmp[267][0][0] = in267;
        tmp[268][0][0] = in268;
        tmp[269][0][0] = in269;
        tmp[270][0][0] = in270;
        tmp[271][0][0] = in271;
        tmp[272][0][0] = in272;
        tmp[273][0][0] = in273;
        tmp[274][0][0] = in274;
        tmp[275][0][0] = in275;
        tmp[276][0][0] = in276;
        tmp[277][0][0] = in277;
        tmp[278][0][0] = in278;
        tmp[279][0][0] = in279;
        tmp[280][0][0] = in280;
        tmp[281][0][0] = in281;
        tmp[282][0][0] = in282;
        tmp[283][0][0] = in283;
        tmp[284][0][0] = in284;
        tmp[285][0][0] = in285;
        tmp[286][0][0] = in286;
        tmp[287][0][0] = in287;
        tmp[288][0][0] = in288;
        tmp[289][0][0] = in289;
        tmp[290][0][0] = in290;
        tmp[291][0][0] = in291;
        tmp[292][0][0] = in292;
        tmp[293][0][0] = in293;
        tmp[294][0][0] = in294;
        tmp[295][0][0] = in295;
        tmp[296][0][0] = in296;
        tmp[297][0][0] = in297;
        tmp[298][0][0] = in298;
        tmp[299][0][0] = in299;
        tmp[300][0][0] = in300;
        tmp[301][0][0] = in301;
        tmp[302][0][0] = in302;
        tmp[303][0][0] = in303;
        tmp[304][0][0] = in304;
        tmp[305][0][0] = in305;
        tmp[306][0][0] = in306;
        tmp[307][0][0] = in307;
        tmp[308][0][0] = in308;
        tmp[309][0][0] = in309;
        tmp[310][0][0] = in310;
        tmp[311][0][0] = in311;
        tmp[312][0][0] = in312;
        tmp[313][0][0] = in313;
        tmp[314][0][0] = in314;
        tmp[315][0][0] = in315;
        tmp[316][0][0] = in316;
        tmp[317][0][0] = in317;
        tmp[318][0][0] = in318;
        tmp[319][0][0] = in319;
        tmp[320][0][0] = in320;
        tmp[321][0][0] = in321;
        tmp[322][0][0] = in322;
        tmp[323][0][0] = in323;
        tmp[324][0][0] = in324;
        tmp[325][0][0] = in325;
        tmp[326][0][0] = in326;
        tmp[327][0][0] = in327;
        tmp[328][0][0] = in328;
        tmp[329][0][0] = in329;
        tmp[330][0][0] = in330;
        tmp[331][0][0] = in331;
        tmp[332][0][0] = in332;
        tmp[333][0][0] = in333;
        tmp[334][0][0] = in334;
        tmp[335][0][0] = in335;
        tmp[336][0][0] = in336;
        tmp[337][0][0] = in337;
        tmp[338][0][0] = in338;
        tmp[339][0][0] = in339;
        tmp[340][0][0] = in340;
        tmp[341][0][0] = in341;
        tmp[342][0][0] = in342;
        tmp[343][0][0] = in343;
        tmp[344][0][0] = in344;
        tmp[345][0][0] = in345;
        tmp[346][0][0] = in346;
        tmp[347][0][0] = in347;
        tmp[348][0][0] = in348;
        tmp[349][0][0] = in349;
        tmp[350][0][0] = in350;
        tmp[351][0][0] = in351;
        tmp[352][0][0] = in352;
        tmp[353][0][0] = in353;
        tmp[354][0][0] = in354;
        tmp[355][0][0] = in355;
        tmp[356][0][0] = in356;
        tmp[357][0][0] = in357;
        tmp[358][0][0] = in358;
        tmp[359][0][0] = in359;
        tmp[360][0][0] = in360;
        tmp[361][0][0] = in361;
        tmp[362][0][0] = in362;
        tmp[363][0][0] = in363;
        tmp[364][0][0] = in364;
        tmp[365][0][0] = in365;
        tmp[366][0][0] = in366;
        tmp[367][0][0] = in367;
        tmp[368][0][0] = in368;
        tmp[369][0][0] = in369;
        tmp[370][0][0] = in370;
        tmp[371][0][0] = in371;
        tmp[372][0][0] = in372;
        tmp[373][0][0] = in373;
        tmp[374][0][0] = in374;
        tmp[375][0][0] = in375;
        tmp[376][0][0] = in376;
        tmp[377][0][0] = in377;
        tmp[378][0][0] = in378;
        tmp[379][0][0] = in379;
        tmp[380][0][0] = in380;
        tmp[381][0][0] = in381;
        tmp[382][0][0] = in382;
        tmp[383][0][0] = in383;
        tmp[384][0][0] = in384;
        tmp[385][0][0] = in385;
        tmp[386][0][0] = in386;
        tmp[387][0][0] = in387;
        tmp[388][0][0] = in388;
        tmp[389][0][0] = in389;
        tmp[390][0][0] = in390;
        tmp[391][0][0] = in391;
        tmp[392][0][0] = in392;
        tmp[393][0][0] = in393;
        tmp[394][0][0] = in394;
        tmp[395][0][0] = in395;
        tmp[396][0][0] = in396;
        tmp[397][0][0] = in397;
        tmp[398][0][0] = in398;
        tmp[399][0][0] = in399;
        tmp[400][0][0] = in400;
        tmp[401][0][0] = in401;
        tmp[402][0][0] = in402;
        tmp[403][0][0] = in403;
        tmp[404][0][0] = in404;
        tmp[405][0][0] = in405;
        tmp[406][0][0] = in406;
        tmp[407][0][0] = in407;
        tmp[408][0][0] = in408;
        tmp[409][0][0] = in409;
        tmp[410][0][0] = in410;
        tmp[411][0][0] = in411;
        tmp[412][0][0] = in412;
        tmp[413][0][0] = in413;
        tmp[414][0][0] = in414;
        tmp[415][0][0] = in415;
        tmp[416][0][0] = in416;
        tmp[417][0][0] = in417;
        tmp[418][0][0] = in418;
        tmp[419][0][0] = in419;
        tmp[420][0][0] = in420;
        tmp[421][0][0] = in421;
        tmp[422][0][0] = in422;
        tmp[423][0][0] = in423;
        tmp[424][0][0] = in424;
        tmp[425][0][0] = in425;
        tmp[426][0][0] = in426;
        tmp[427][0][0] = in427;
        tmp[428][0][0] = in428;
        tmp[429][0][0] = in429;
        tmp[430][0][0] = in430;
        tmp[431][0][0] = in431;
        tmp[432][0][0] = in432;
        tmp[433][0][0] = in433;
        tmp[434][0][0] = in434;
        tmp[435][0][0] = in435;
        tmp[436][0][0] = in436;
        tmp[437][0][0] = in437;
        tmp[438][0][0] = in438;
        tmp[439][0][0] = in439;
        tmp[440][0][0] = in440;
        tmp[441][0][0] = in441;
        tmp[442][0][0] = in442;
        tmp[443][0][0] = in443;
        tmp[444][0][0] = in444;
        tmp[445][0][0] = in445;
        tmp[446][0][0] = in446;
        tmp[447][0][0] = in447;
        tmp[448][0][0] = in448;
        tmp[449][0][0] = in449;
        tmp[450][0][0] = in450;
        tmp[451][0][0] = in451;
        tmp[452][0][0] = in452;
        tmp[453][0][0] = in453;
        tmp[454][0][0] = in454;
        tmp[455][0][0] = in455;
        tmp[456][0][0] = in456;
        tmp[457][0][0] = in457;
        tmp[458][0][0] = in458;
        tmp[459][0][0] = in459;
        tmp[460][0][0] = in460;
        tmp[461][0][0] = in461;
        tmp[462][0][0] = in462;
        tmp[463][0][0] = in463;
        tmp[464][0][0] = in464;
        tmp[465][0][0] = in465;
        tmp[466][0][0] = in466;
        tmp[467][0][0] = in467;
        tmp[468][0][0] = in468;
        tmp[469][0][0] = in469;
        tmp[470][0][0] = in470;
        tmp[471][0][0] = in471;
        tmp[472][0][0] = in472;
        tmp[473][0][0] = in473;
        tmp[474][0][0] = in474;
        tmp[475][0][0] = in475;
        tmp[476][0][0] = in476;
        tmp[477][0][0] = in477;
        tmp[478][0][0] = in478;
        tmp[479][0][0] = in479;
        tmp[480][0][0] = in480;
        tmp[481][0][0] = in481;
        tmp[482][0][0] = in482;
        tmp[483][0][0] = in483;
        tmp[484][0][0] = in484;
        tmp[485][0][0] = in485;
        tmp[486][0][0] = in486;
        tmp[487][0][0] = in487;
        tmp[488][0][0] = in488;
        tmp[489][0][0] = in489;
        tmp[490][0][0] = in490;
        tmp[491][0][0] = in491;
        tmp[492][0][0] = in492;
        tmp[493][0][0] = in493;
        tmp[494][0][0] = in494;
        tmp[495][0][0] = in495;
        tmp[496][0][0] = in496;
        tmp[497][0][0] = in497;
        tmp[498][0][0] = in498;
        tmp[499][0][0] = in499;
        tmp[500][0][0] = in500;
        tmp[501][0][0] = in501;
        tmp[502][0][0] = in502;
        tmp[503][0][0] = in503;
        tmp[504][0][0] = in504;
        tmp[505][0][0] = in505;
        tmp[506][0][0] = in506;
        tmp[507][0][0] = in507;
        tmp[508][0][0] = in508;
        tmp[509][0][0] = in509;
        tmp[510][0][0] = in510;
        tmp[511][0][0] = in511;
        tmp[512][0][0] = in512;
        tmp[513][0][0] = in513;
        tmp[514][0][0] = in514;
        tmp[515][0][0] = in515;
        tmp[516][0][0] = in516;
        tmp[517][0][0] = in517;
        tmp[518][0][0] = in518;
        tmp[519][0][0] = in519;
        tmp[520][0][0] = in520;
        tmp[521][0][0] = in521;
        tmp[522][0][0] = in522;
        tmp[523][0][0] = in523;
        tmp[524][0][0] = in524;
        tmp[525][0][0] = in525;
        tmp[526][0][0] = in526;
        tmp[527][0][0] = in527;
        tmp[528][0][0] = in528;
        tmp[529][0][0] = in529;
        tmp[530][0][0] = in530;
        tmp[531][0][0] = in531;
        tmp[532][0][0] = in532;
        tmp[533][0][0] = in533;
        tmp[534][0][0] = in534;
        tmp[535][0][0] = in535;
        tmp[536][0][0] = in536;
        tmp[537][0][0] = in537;
        tmp[538][0][0] = in538;
        tmp[539][0][0] = in539;
        tmp[540][0][0] = in540;
        tmp[541][0][0] = in541;
        tmp[542][0][0] = in542;
        tmp[543][0][0] = in543;
        tmp[544][0][0] = in544;
        tmp[545][0][0] = in545;
        tmp[546][0][0] = in546;
        tmp[547][0][0] = in547;
        tmp[548][0][0] = in548;
        tmp[549][0][0] = in549;
        tmp[550][0][0] = in550;
        tmp[551][0][0] = in551;
        tmp[552][0][0] = in552;
        tmp[553][0][0] = in553;
        tmp[554][0][0] = in554;
        tmp[555][0][0] = in555;
        tmp[556][0][0] = in556;
        tmp[557][0][0] = in557;
        tmp[558][0][0] = in558;
        tmp[559][0][0] = in559;
        tmp[560][0][0] = in560;
        tmp[561][0][0] = in561;
        tmp[562][0][0] = in562;
        tmp[563][0][0] = in563;
        tmp[564][0][0] = in564;
        tmp[565][0][0] = in565;
        tmp[566][0][0] = in566;
        tmp[567][0][0] = in567;
        tmp[568][0][0] = in568;
        tmp[569][0][0] = in569;
        tmp[570][0][0] = in570;
        tmp[571][0][0] = in571;
        tmp[572][0][0] = in572;
        tmp[573][0][0] = in573;
        tmp[574][0][0] = in574;
        tmp[575][0][0] = in575;
        tmp[576][0][0] = in576;
        tmp[577][0][0] = in577;
        tmp[578][0][0] = in578;
        tmp[579][0][0] = in579;
        tmp[580][0][0] = in580;
        tmp[581][0][0] = in581;
        tmp[582][0][0] = in582;
        tmp[583][0][0] = in583;
        tmp[584][0][0] = in584;
        tmp[585][0][0] = in585;
        tmp[586][0][0] = in586;
        tmp[587][0][0] = in587;
        tmp[588][0][0] = in588;
        tmp[589][0][0] = in589;
        tmp[590][0][0] = in590;
        tmp[591][0][0] = in591;
        tmp[592][0][0] = in592;
        tmp[593][0][0] = in593;
        tmp[594][0][0] = in594;
        tmp[595][0][0] = in595;
        tmp[596][0][0] = in596;
        tmp[597][0][0] = in597;
        tmp[598][0][0] = in598;
        tmp[599][0][0] = in599;
        tmp[600][0][0] = in600;
        tmp[601][0][0] = in601;
        tmp[602][0][0] = in602;
        tmp[603][0][0] = in603;
        tmp[604][0][0] = in604;
        tmp[605][0][0] = in605;
        tmp[606][0][0] = in606;
        tmp[607][0][0] = in607;
        tmp[608][0][0] = in608;
        tmp[609][0][0] = in609;
        tmp[610][0][0] = in610;
        tmp[611][0][0] = in611;
        tmp[612][0][0] = in612;
        tmp[613][0][0] = in613;
        tmp[614][0][0] = in614;
        tmp[615][0][0] = in615;
        tmp[616][0][0] = in616;
        tmp[617][0][0] = in617;
        tmp[618][0][0] = in618;
        tmp[619][0][0] = in619;
        tmp[620][0][0] = in620;
        tmp[621][0][0] = in621;
        tmp[622][0][0] = in622;
        tmp[623][0][0] = in623;
        tmp[624][0][0] = in624;
        tmp[625][0][0] = in625;
        tmp[626][0][0] = in626;
        tmp[627][0][0] = in627;
        tmp[628][0][0] = in628;
        tmp[629][0][0] = in629;
        tmp[630][0][0] = in630;
        tmp[631][0][0] = in631;
        tmp[632][0][0] = in632;
        tmp[633][0][0] = in633;
        tmp[634][0][0] = in634;
        tmp[635][0][0] = in635;
        tmp[636][0][0] = in636;
        tmp[637][0][0] = in637;
        tmp[638][0][0] = in638;
        tmp[639][0][0] = in639;
        tmp[640][0][0] = in640;
        tmp[641][0][0] = in641;
        tmp[642][0][0] = in642;
        tmp[643][0][0] = in643;
        tmp[644][0][0] = in644;
        tmp[645][0][0] = in645;
        tmp[646][0][0] = in646;
        tmp[647][0][0] = in647;
        tmp[648][0][0] = in648;
        tmp[649][0][0] = in649;
        tmp[650][0][0] = in650;
        tmp[651][0][0] = in651;
        tmp[652][0][0] = in652;
        tmp[653][0][0] = in653;
        tmp[654][0][0] = in654;
        tmp[655][0][0] = in655;
        tmp[656][0][0] = in656;
        tmp[657][0][0] = in657;
        tmp[658][0][0] = in658;
        tmp[659][0][0] = in659;
        tmp[660][0][0] = in660;
        tmp[661][0][0] = in661;
        tmp[662][0][0] = in662;
        tmp[663][0][0] = in663;
        tmp[664][0][0] = in664;
        tmp[665][0][0] = in665;
        tmp[666][0][0] = in666;
        tmp[667][0][0] = in667;
        tmp[668][0][0] = in668;
        tmp[669][0][0] = in669;
        tmp[670][0][0] = in670;
        tmp[671][0][0] = in671;
        tmp[672][0][0] = in672;
        tmp[673][0][0] = in673;
        tmp[674][0][0] = in674;
        tmp[675][0][0] = in675;
        tmp[676][0][0] = in676;
        tmp[677][0][0] = in677;
        tmp[678][0][0] = in678;
        tmp[679][0][0] = in679;
        tmp[680][0][0] = in680;
        tmp[681][0][0] = in681;
        tmp[682][0][0] = in682;
        tmp[683][0][0] = in683;
        tmp[684][0][0] = in684;
        tmp[685][0][0] = in685;
        tmp[686][0][0] = in686;
        tmp[687][0][0] = in687;
        tmp[688][0][0] = in688;
        tmp[689][0][0] = in689;
        tmp[690][0][0] = in690;
        tmp[691][0][0] = in691;
        tmp[692][0][0] = in692;
        tmp[693][0][0] = in693;
        tmp[694][0][0] = in694;
        tmp[695][0][0] = in695;
        tmp[696][0][0] = in696;
        tmp[697][0][0] = in697;
        tmp[698][0][0] = in698;
        tmp[699][0][0] = in699;
        tmp[700][0][0] = in700;
        tmp[701][0][0] = in701;
        tmp[702][0][0] = in702;
        tmp[703][0][0] = in703;
        tmp[704][0][0] = in704;
        tmp[705][0][0] = in705;
        tmp[706][0][0] = in706;
        tmp[707][0][0] = in707;
        tmp[708][0][0] = in708;
        tmp[709][0][0] = in709;
        tmp[710][0][0] = in710;
        tmp[711][0][0] = in711;
        tmp[712][0][0] = in712;
        tmp[713][0][0] = in713;
        tmp[714][0][0] = in714;
        tmp[715][0][0] = in715;
        tmp[716][0][0] = in716;
        tmp[717][0][0] = in717;
        tmp[718][0][0] = in718;
        tmp[719][0][0] = in719;
        tmp[720][0][0] = in720;
        tmp[721][0][0] = in721;
        tmp[722][0][0] = in722;
        tmp[723][0][0] = in723;
        tmp[724][0][0] = in724;
        tmp[725][0][0] = in725;
        tmp[726][0][0] = in726;
        tmp[727][0][0] = in727;
        tmp[728][0][0] = in728;
        tmp[729][0][0] = in729;
        tmp[730][0][0] = in730;
        tmp[731][0][0] = in731;
        tmp[732][0][0] = in732;
        tmp[733][0][0] = in733;
        tmp[734][0][0] = in734;
        tmp[735][0][0] = in735;
        tmp[736][0][0] = in736;
        tmp[737][0][0] = in737;
        tmp[738][0][0] = in738;
        tmp[739][0][0] = in739;
        tmp[740][0][0] = in740;
        tmp[741][0][0] = in741;
        tmp[742][0][0] = in742;
        tmp[743][0][0] = in743;
        tmp[744][0][0] = in744;
        tmp[745][0][0] = in745;
        tmp[746][0][0] = in746;
        tmp[747][0][0] = in747;
        tmp[748][0][0] = in748;
        tmp[749][0][0] = in749;
        tmp[750][0][0] = in750;
        tmp[751][0][0] = in751;
        tmp[752][0][0] = in752;
        tmp[753][0][0] = in753;
        tmp[754][0][0] = in754;
        tmp[755][0][0] = in755;
        tmp[756][0][0] = in756;
        tmp[757][0][0] = in757;
        tmp[758][0][0] = in758;
        tmp[759][0][0] = in759;
        tmp[760][0][0] = in760;
        tmp[761][0][0] = in761;
        tmp[762][0][0] = in762;
        tmp[763][0][0] = in763;
        tmp[764][0][0] = in764;
        tmp[765][0][0] = in765;
        tmp[766][0][0] = in766;
        tmp[767][0][0] = in767;
        tmp[768][0][0] = in768;
        tmp[769][0][0] = in769;
        tmp[770][0][0] = in770;
        tmp[771][0][0] = in771;
        tmp[772][0][0] = in772;
        tmp[773][0][0] = in773;
        tmp[774][0][0] = in774;
        tmp[775][0][0] = in775;
        tmp[776][0][0] = in776;
        tmp[777][0][0] = in777;
        tmp[778][0][0] = in778;
        tmp[779][0][0] = in779;
        tmp[780][0][0] = in780;
        tmp[781][0][0] = in781;
        tmp[782][0][0] = in782;
        tmp[783][0][0] = in783;
        tmp[784][0][0] = in784;
        tmp[785][0][0] = in785;
        tmp[786][0][0] = in786;
        tmp[787][0][0] = in787;
        tmp[788][0][0] = in788;
        tmp[789][0][0] = in789;
        tmp[790][0][0] = in790;
        tmp[791][0][0] = in791;
        tmp[792][0][0] = in792;
        tmp[793][0][0] = in793;
        tmp[794][0][0] = in794;
        tmp[795][0][0] = in795;
        tmp[796][0][0] = in796;
        tmp[797][0][0] = in797;
        tmp[798][0][0] = in798;
        tmp[799][0][0] = in799;
        tmp[800][0][0] = in800;
        tmp[801][0][0] = in801;
        tmp[802][0][0] = in802;
        tmp[803][0][0] = in803;
        tmp[804][0][0] = in804;
        tmp[805][0][0] = in805;
        tmp[806][0][0] = in806;
        tmp[807][0][0] = in807;
        tmp[808][0][0] = in808;
        tmp[809][0][0] = in809;
        tmp[810][0][0] = in810;
        tmp[811][0][0] = in811;
        tmp[812][0][0] = in812;
        tmp[813][0][0] = in813;
        tmp[814][0][0] = in814;
        tmp[815][0][0] = in815;
        tmp[816][0][0] = in816;
        tmp[817][0][0] = in817;
        tmp[818][0][0] = in818;
        tmp[819][0][0] = in819;
        tmp[820][0][0] = in820;
        tmp[821][0][0] = in821;
        tmp[822][0][0] = in822;
        tmp[823][0][0] = in823;
        tmp[824][0][0] = in824;
        tmp[825][0][0] = in825;
        tmp[826][0][0] = in826;
        tmp[827][0][0] = in827;
        tmp[828][0][0] = in828;
        tmp[829][0][0] = in829;
        tmp[830][0][0] = in830;
        tmp[831][0][0] = in831;
        tmp[832][0][0] = in832;
        tmp[833][0][0] = in833;
        tmp[834][0][0] = in834;
        tmp[835][0][0] = in835;
        tmp[836][0][0] = in836;
        tmp[837][0][0] = in837;
        tmp[838][0][0] = in838;
        tmp[839][0][0] = in839;
        tmp[840][0][0] = in840;
        tmp[841][0][0] = in841;
        tmp[842][0][0] = in842;
        tmp[843][0][0] = in843;
        tmp[844][0][0] = in844;
        tmp[845][0][0] = in845;
        tmp[846][0][0] = in846;
        tmp[847][0][0] = in847;
        tmp[848][0][0] = in848;
        tmp[849][0][0] = in849;
        tmp[850][0][0] = in850;
        tmp[851][0][0] = in851;
        tmp[852][0][0] = in852;
        tmp[853][0][0] = in853;
        tmp[854][0][0] = in854;
        tmp[855][0][0] = in855;
        tmp[856][0][0] = in856;
        tmp[857][0][0] = in857;
        tmp[858][0][0] = in858;
        tmp[859][0][0] = in859;
        tmp[860][0][0] = in860;
        tmp[861][0][0] = in861;
        tmp[862][0][0] = in862;
        tmp[863][0][0] = in863;
        tmp[864][0][0] = in864;
        tmp[865][0][0] = in865;
        tmp[866][0][0] = in866;
        tmp[867][0][0] = in867;
        tmp[868][0][0] = in868;
        tmp[869][0][0] = in869;
        tmp[870][0][0] = in870;
        tmp[871][0][0] = in871;
        tmp[872][0][0] = in872;
        tmp[873][0][0] = in873;
        tmp[874][0][0] = in874;
        tmp[875][0][0] = in875;
        tmp[876][0][0] = in876;
        tmp[877][0][0] = in877;
        tmp[878][0][0] = in878;
        tmp[879][0][0] = in879;
        tmp[880][0][0] = in880;
        tmp[881][0][0] = in881;
        tmp[882][0][0] = in882;
        tmp[883][0][0] = in883;
        tmp[884][0][0] = in884;
        tmp[885][0][0] = in885;
        tmp[886][0][0] = in886;
        tmp[887][0][0] = in887;
        tmp[888][0][0] = in888;
        tmp[889][0][0] = in889;
        tmp[890][0][0] = in890;
        tmp[891][0][0] = in891;
        tmp[892][0][0] = in892;
        tmp[893][0][0] = in893;
        tmp[894][0][0] = in894;
        tmp[895][0][0] = in895;
        tmp[896][0][0] = in896;
        tmp[897][0][0] = in897;
        tmp[898][0][0] = in898;
        tmp[899][0][0] = in899;
        tmp[900][0][0] = in900;
        tmp[901][0][0] = in901;
        tmp[902][0][0] = in902;
        tmp[903][0][0] = in903;
        tmp[904][0][0] = in904;
        tmp[905][0][0] = in905;
        tmp[906][0][0] = in906;
        tmp[907][0][0] = in907;
        tmp[908][0][0] = in908;
        tmp[909][0][0] = in909;
        tmp[910][0][0] = in910;
        tmp[911][0][0] = in911;
        tmp[912][0][0] = in912;
        tmp[913][0][0] = in913;
        tmp[914][0][0] = in914;
        tmp[915][0][0] = in915;
        tmp[916][0][0] = in916;
        tmp[917][0][0] = in917;
        tmp[918][0][0] = in918;
        tmp[919][0][0] = in919;
        tmp[920][0][0] = in920;
        tmp[921][0][0] = in921;
        tmp[922][0][0] = in922;
        tmp[923][0][0] = in923;
        tmp[924][0][0] = in924;
        tmp[925][0][0] = in925;
        tmp[926][0][0] = in926;
        tmp[927][0][0] = in927;
        tmp[928][0][0] = in928;
        tmp[929][0][0] = in929;
        tmp[930][0][0] = in930;
        tmp[931][0][0] = in931;
        tmp[932][0][0] = in932;
        tmp[933][0][0] = in933;
        tmp[934][0][0] = in934;
        tmp[935][0][0] = in935;
        tmp[936][0][0] = in936;
        tmp[937][0][0] = in937;
        tmp[938][0][0] = in938;
        tmp[939][0][0] = in939;
        tmp[940][0][0] = in940;
        tmp[941][0][0] = in941;
        tmp[942][0][0] = in942;
        tmp[943][0][0] = in943;
        tmp[944][0][0] = in944;
        tmp[945][0][0] = in945;
        tmp[946][0][0] = in946;
        tmp[947][0][0] = in947;
        tmp[948][0][0] = in948;
        tmp[949][0][0] = in949;
        tmp[950][0][0] = in950;
        tmp[951][0][0] = in951;
        tmp[952][0][0] = in952;
        tmp[953][0][0] = in953;
        tmp[954][0][0] = in954;
        tmp[955][0][0] = in955;
        tmp[956][0][0] = in956;
        tmp[957][0][0] = in957;
        tmp[958][0][0] = in958;
        tmp[959][0][0] = in959;
        tmp[960][0][0] = in960;
        tmp[961][0][0] = in961;
        tmp[962][0][0] = in962;
        tmp[963][0][0] = in963;
        tmp[964][0][0] = in964;
        tmp[965][0][0] = in965;
        tmp[966][0][0] = in966;
        tmp[967][0][0] = in967;
        tmp[968][0][0] = in968;
        tmp[969][0][0] = in969;
        tmp[970][0][0] = in970;
        tmp[971][0][0] = in971;
        tmp[972][0][0] = in972;
        tmp[973][0][0] = in973;
        tmp[974][0][0] = in974;
        tmp[975][0][0] = in975;
        tmp[976][0][0] = in976;
        tmp[977][0][0] = in977;
        tmp[978][0][0] = in978;
        tmp[979][0][0] = in979;
        tmp[980][0][0] = in980;
        tmp[981][0][0] = in981;
        tmp[982][0][0] = in982;
        tmp[983][0][0] = in983;
        tmp[984][0][0] = in984;
        tmp[985][0][0] = in985;
        tmp[986][0][0] = in986;
        tmp[987][0][0] = in987;
        tmp[988][0][0] = in988;
        tmp[989][0][0] = in989;
        tmp[990][0][0] = in990;
        tmp[991][0][0] = in991;
        tmp[992][0][0] = in992;
        tmp[993][0][0] = in993;
        tmp[994][0][0] = in994;
        tmp[995][0][0] = in995;
        tmp[996][0][0] = in996;
        tmp[997][0][0] = in997;
        tmp[998][0][0] = in998;
        tmp[999][0][0] = in999;
        tmp[1000][0][0] = in1000;
        tmp[1001][0][0] = in1001;
        tmp[1002][0][0] = in1002;
        tmp[1003][0][0] = in1003;
        tmp[1004][0][0] = in1004;
        tmp[1005][0][0] = in1005;
        tmp[1006][0][0] = in1006;
        tmp[1007][0][0] = in1007;
        tmp[1008][0][0] = in1008;
        tmp[1009][0][0] = in1009;
        tmp[1010][0][0] = in1010;
        tmp[1011][0][0] = in1011;
        tmp[1012][0][0] = in1012;
        tmp[1013][0][0] = in1013;
        tmp[1014][0][0] = in1014;
        tmp[1015][0][0] = in1015;
        tmp[1016][0][0] = in1016;
        tmp[1017][0][0] = in1017;
        tmp[1018][0][0] = in1018;
        tmp[1019][0][0] = in1019;
        tmp[1020][0][0] = in1020;
        tmp[1021][0][0] = in1021;
        tmp[1022][0][0] = in1022;
        tmp[1023][0][0] = in1023;
    end
    assign out0 = tmp[0][STEP][0];
    assign out1 = tmp[1][STEP][0];
    assign out2 = tmp[2][STEP][0];
    assign out3 = tmp[3][STEP][0];
    assign out4 = tmp[4][STEP][0];
    assign out5 = tmp[5][STEP][0];
    assign out6 = tmp[6][STEP][0];
    assign out7 = tmp[7][STEP][0];
    assign out8 = tmp[8][STEP][0];
    assign out9 = tmp[9][STEP][0];
    assign out10 = tmp[10][STEP][0];
    assign out11 = tmp[11][STEP][0];
    assign out12 = tmp[12][STEP][0];
    assign out13 = tmp[13][STEP][0];
    assign out14 = tmp[14][STEP][0];
    assign out15 = tmp[15][STEP][0];
    assign out16 = tmp[16][STEP][0];
    assign out17 = tmp[17][STEP][0];
    assign out18 = tmp[18][STEP][0];
    assign out19 = tmp[19][STEP][0];
    assign out20 = tmp[20][STEP][0];
    assign out21 = tmp[21][STEP][0];
    assign out22 = tmp[22][STEP][0];
    assign out23 = tmp[23][STEP][0];
    assign out24 = tmp[24][STEP][0];
    assign out25 = tmp[25][STEP][0];
    assign out26 = tmp[26][STEP][0];
    assign out27 = tmp[27][STEP][0];
    assign out28 = tmp[28][STEP][0];
    assign out29 = tmp[29][STEP][0];
    assign out30 = tmp[30][STEP][0];
    assign out31 = tmp[31][STEP][0];
    assign out32 = tmp[32][STEP][0];
    assign out33 = tmp[33][STEP][0];
    assign out34 = tmp[34][STEP][0];
    assign out35 = tmp[35][STEP][0];
    assign out36 = tmp[36][STEP][0];
    assign out37 = tmp[37][STEP][0];
    assign out38 = tmp[38][STEP][0];
    assign out39 = tmp[39][STEP][0];
    assign out40 = tmp[40][STEP][0];
    assign out41 = tmp[41][STEP][0];
    assign out42 = tmp[42][STEP][0];
    assign out43 = tmp[43][STEP][0];
    assign out44 = tmp[44][STEP][0];
    assign out45 = tmp[45][STEP][0];
    assign out46 = tmp[46][STEP][0];
    assign out47 = tmp[47][STEP][0];
    assign out48 = tmp[48][STEP][0];
    assign out49 = tmp[49][STEP][0];
    assign out50 = tmp[50][STEP][0];
    assign out51 = tmp[51][STEP][0];
    assign out52 = tmp[52][STEP][0];
    assign out53 = tmp[53][STEP][0];
    assign out54 = tmp[54][STEP][0];
    assign out55 = tmp[55][STEP][0];
    assign out56 = tmp[56][STEP][0];
    assign out57 = tmp[57][STEP][0];
    assign out58 = tmp[58][STEP][0];
    assign out59 = tmp[59][STEP][0];
    assign out60 = tmp[60][STEP][0];
    assign out61 = tmp[61][STEP][0];
    assign out62 = tmp[62][STEP][0];
    assign out63 = tmp[63][STEP][0];
    assign out64 = tmp[64][STEP][0];
    assign out65 = tmp[65][STEP][0];
    assign out66 = tmp[66][STEP][0];
    assign out67 = tmp[67][STEP][0];
    assign out68 = tmp[68][STEP][0];
    assign out69 = tmp[69][STEP][0];
    assign out70 = tmp[70][STEP][0];
    assign out71 = tmp[71][STEP][0];
    assign out72 = tmp[72][STEP][0];
    assign out73 = tmp[73][STEP][0];
    assign out74 = tmp[74][STEP][0];
    assign out75 = tmp[75][STEP][0];
    assign out76 = tmp[76][STEP][0];
    assign out77 = tmp[77][STEP][0];
    assign out78 = tmp[78][STEP][0];
    assign out79 = tmp[79][STEP][0];
    assign out80 = tmp[80][STEP][0];
    assign out81 = tmp[81][STEP][0];
    assign out82 = tmp[82][STEP][0];
    assign out83 = tmp[83][STEP][0];
    assign out84 = tmp[84][STEP][0];
    assign out85 = tmp[85][STEP][0];
    assign out86 = tmp[86][STEP][0];
    assign out87 = tmp[87][STEP][0];
    assign out88 = tmp[88][STEP][0];
    assign out89 = tmp[89][STEP][0];
    assign out90 = tmp[90][STEP][0];
    assign out91 = tmp[91][STEP][0];
    assign out92 = tmp[92][STEP][0];
    assign out93 = tmp[93][STEP][0];
    assign out94 = tmp[94][STEP][0];
    assign out95 = tmp[95][STEP][0];
    assign out96 = tmp[96][STEP][0];
    assign out97 = tmp[97][STEP][0];
    assign out98 = tmp[98][STEP][0];
    assign out99 = tmp[99][STEP][0];
    assign out100 = tmp[100][STEP][0];
    assign out101 = tmp[101][STEP][0];
    assign out102 = tmp[102][STEP][0];
    assign out103 = tmp[103][STEP][0];
    assign out104 = tmp[104][STEP][0];
    assign out105 = tmp[105][STEP][0];
    assign out106 = tmp[106][STEP][0];
    assign out107 = tmp[107][STEP][0];
    assign out108 = tmp[108][STEP][0];
    assign out109 = tmp[109][STEP][0];
    assign out110 = tmp[110][STEP][0];
    assign out111 = tmp[111][STEP][0];
    assign out112 = tmp[112][STEP][0];
    assign out113 = tmp[113][STEP][0];
    assign out114 = tmp[114][STEP][0];
    assign out115 = tmp[115][STEP][0];
    assign out116 = tmp[116][STEP][0];
    assign out117 = tmp[117][STEP][0];
    assign out118 = tmp[118][STEP][0];
    assign out119 = tmp[119][STEP][0];
    assign out120 = tmp[120][STEP][0];
    assign out121 = tmp[121][STEP][0];
    assign out122 = tmp[122][STEP][0];
    assign out123 = tmp[123][STEP][0];
    assign out124 = tmp[124][STEP][0];
    assign out125 = tmp[125][STEP][0];
    assign out126 = tmp[126][STEP][0];
    assign out127 = tmp[127][STEP][0];
    assign out128 = tmp[128][STEP][0];
    assign out129 = tmp[129][STEP][0];
    assign out130 = tmp[130][STEP][0];
    assign out131 = tmp[131][STEP][0];
    assign out132 = tmp[132][STEP][0];
    assign out133 = tmp[133][STEP][0];
    assign out134 = tmp[134][STEP][0];
    assign out135 = tmp[135][STEP][0];
    assign out136 = tmp[136][STEP][0];
    assign out137 = tmp[137][STEP][0];
    assign out138 = tmp[138][STEP][0];
    assign out139 = tmp[139][STEP][0];
    assign out140 = tmp[140][STEP][0];
    assign out141 = tmp[141][STEP][0];
    assign out142 = tmp[142][STEP][0];
    assign out143 = tmp[143][STEP][0];
    assign out144 = tmp[144][STEP][0];
    assign out145 = tmp[145][STEP][0];
    assign out146 = tmp[146][STEP][0];
    assign out147 = tmp[147][STEP][0];
    assign out148 = tmp[148][STEP][0];
    assign out149 = tmp[149][STEP][0];
    assign out150 = tmp[150][STEP][0];
    assign out151 = tmp[151][STEP][0];
    assign out152 = tmp[152][STEP][0];
    assign out153 = tmp[153][STEP][0];
    assign out154 = tmp[154][STEP][0];
    assign out155 = tmp[155][STEP][0];
    assign out156 = tmp[156][STEP][0];
    assign out157 = tmp[157][STEP][0];
    assign out158 = tmp[158][STEP][0];
    assign out159 = tmp[159][STEP][0];
    assign out160 = tmp[160][STEP][0];
    assign out161 = tmp[161][STEP][0];
    assign out162 = tmp[162][STEP][0];
    assign out163 = tmp[163][STEP][0];
    assign out164 = tmp[164][STEP][0];
    assign out165 = tmp[165][STEP][0];
    assign out166 = tmp[166][STEP][0];
    assign out167 = tmp[167][STEP][0];
    assign out168 = tmp[168][STEP][0];
    assign out169 = tmp[169][STEP][0];
    assign out170 = tmp[170][STEP][0];
    assign out171 = tmp[171][STEP][0];
    assign out172 = tmp[172][STEP][0];
    assign out173 = tmp[173][STEP][0];
    assign out174 = tmp[174][STEP][0];
    assign out175 = tmp[175][STEP][0];
    assign out176 = tmp[176][STEP][0];
    assign out177 = tmp[177][STEP][0];
    assign out178 = tmp[178][STEP][0];
    assign out179 = tmp[179][STEP][0];
    assign out180 = tmp[180][STEP][0];
    assign out181 = tmp[181][STEP][0];
    assign out182 = tmp[182][STEP][0];
    assign out183 = tmp[183][STEP][0];
    assign out184 = tmp[184][STEP][0];
    assign out185 = tmp[185][STEP][0];
    assign out186 = tmp[186][STEP][0];
    assign out187 = tmp[187][STEP][0];
    assign out188 = tmp[188][STEP][0];
    assign out189 = tmp[189][STEP][0];
    assign out190 = tmp[190][STEP][0];
    assign out191 = tmp[191][STEP][0];
    assign out192 = tmp[192][STEP][0];
    assign out193 = tmp[193][STEP][0];
    assign out194 = tmp[194][STEP][0];
    assign out195 = tmp[195][STEP][0];
    assign out196 = tmp[196][STEP][0];
    assign out197 = tmp[197][STEP][0];
    assign out198 = tmp[198][STEP][0];
    assign out199 = tmp[199][STEP][0];
    assign out200 = tmp[200][STEP][0];
    assign out201 = tmp[201][STEP][0];
    assign out202 = tmp[202][STEP][0];
    assign out203 = tmp[203][STEP][0];
    assign out204 = tmp[204][STEP][0];
    assign out205 = tmp[205][STEP][0];
    assign out206 = tmp[206][STEP][0];
    assign out207 = tmp[207][STEP][0];
    assign out208 = tmp[208][STEP][0];
    assign out209 = tmp[209][STEP][0];
    assign out210 = tmp[210][STEP][0];
    assign out211 = tmp[211][STEP][0];
    assign out212 = tmp[212][STEP][0];
    assign out213 = tmp[213][STEP][0];
    assign out214 = tmp[214][STEP][0];
    assign out215 = tmp[215][STEP][0];
    assign out216 = tmp[216][STEP][0];
    assign out217 = tmp[217][STEP][0];
    assign out218 = tmp[218][STEP][0];
    assign out219 = tmp[219][STEP][0];
    assign out220 = tmp[220][STEP][0];
    assign out221 = tmp[221][STEP][0];
    assign out222 = tmp[222][STEP][0];
    assign out223 = tmp[223][STEP][0];
    assign out224 = tmp[224][STEP][0];
    assign out225 = tmp[225][STEP][0];
    assign out226 = tmp[226][STEP][0];
    assign out227 = tmp[227][STEP][0];
    assign out228 = tmp[228][STEP][0];
    assign out229 = tmp[229][STEP][0];
    assign out230 = tmp[230][STEP][0];
    assign out231 = tmp[231][STEP][0];
    assign out232 = tmp[232][STEP][0];
    assign out233 = tmp[233][STEP][0];
    assign out234 = tmp[234][STEP][0];
    assign out235 = tmp[235][STEP][0];
    assign out236 = tmp[236][STEP][0];
    assign out237 = tmp[237][STEP][0];
    assign out238 = tmp[238][STEP][0];
    assign out239 = tmp[239][STEP][0];
    assign out240 = tmp[240][STEP][0];
    assign out241 = tmp[241][STEP][0];
    assign out242 = tmp[242][STEP][0];
    assign out243 = tmp[243][STEP][0];
    assign out244 = tmp[244][STEP][0];
    assign out245 = tmp[245][STEP][0];
    assign out246 = tmp[246][STEP][0];
    assign out247 = tmp[247][STEP][0];
    assign out248 = tmp[248][STEP][0];
    assign out249 = tmp[249][STEP][0];
    assign out250 = tmp[250][STEP][0];
    assign out251 = tmp[251][STEP][0];
    assign out252 = tmp[252][STEP][0];
    assign out253 = tmp[253][STEP][0];
    assign out254 = tmp[254][STEP][0];
    assign out255 = tmp[255][STEP][0];
    assign out256 = tmp[256][STEP][0];
    assign out257 = tmp[257][STEP][0];
    assign out258 = tmp[258][STEP][0];
    assign out259 = tmp[259][STEP][0];
    assign out260 = tmp[260][STEP][0];
    assign out261 = tmp[261][STEP][0];
    assign out262 = tmp[262][STEP][0];
    assign out263 = tmp[263][STEP][0];
    assign out264 = tmp[264][STEP][0];
    assign out265 = tmp[265][STEP][0];
    assign out266 = tmp[266][STEP][0];
    assign out267 = tmp[267][STEP][0];
    assign out268 = tmp[268][STEP][0];
    assign out269 = tmp[269][STEP][0];
    assign out270 = tmp[270][STEP][0];
    assign out271 = tmp[271][STEP][0];
    assign out272 = tmp[272][STEP][0];
    assign out273 = tmp[273][STEP][0];
    assign out274 = tmp[274][STEP][0];
    assign out275 = tmp[275][STEP][0];
    assign out276 = tmp[276][STEP][0];
    assign out277 = tmp[277][STEP][0];
    assign out278 = tmp[278][STEP][0];
    assign out279 = tmp[279][STEP][0];
    assign out280 = tmp[280][STEP][0];
    assign out281 = tmp[281][STEP][0];
    assign out282 = tmp[282][STEP][0];
    assign out283 = tmp[283][STEP][0];
    assign out284 = tmp[284][STEP][0];
    assign out285 = tmp[285][STEP][0];
    assign out286 = tmp[286][STEP][0];
    assign out287 = tmp[287][STEP][0];
    assign out288 = tmp[288][STEP][0];
    assign out289 = tmp[289][STEP][0];
    assign out290 = tmp[290][STEP][0];
    assign out291 = tmp[291][STEP][0];
    assign out292 = tmp[292][STEP][0];
    assign out293 = tmp[293][STEP][0];
    assign out294 = tmp[294][STEP][0];
    assign out295 = tmp[295][STEP][0];
    assign out296 = tmp[296][STEP][0];
    assign out297 = tmp[297][STEP][0];
    assign out298 = tmp[298][STEP][0];
    assign out299 = tmp[299][STEP][0];
    assign out300 = tmp[300][STEP][0];
    assign out301 = tmp[301][STEP][0];
    assign out302 = tmp[302][STEP][0];
    assign out303 = tmp[303][STEP][0];
    assign out304 = tmp[304][STEP][0];
    assign out305 = tmp[305][STEP][0];
    assign out306 = tmp[306][STEP][0];
    assign out307 = tmp[307][STEP][0];
    assign out308 = tmp[308][STEP][0];
    assign out309 = tmp[309][STEP][0];
    assign out310 = tmp[310][STEP][0];
    assign out311 = tmp[311][STEP][0];
    assign out312 = tmp[312][STEP][0];
    assign out313 = tmp[313][STEP][0];
    assign out314 = tmp[314][STEP][0];
    assign out315 = tmp[315][STEP][0];
    assign out316 = tmp[316][STEP][0];
    assign out317 = tmp[317][STEP][0];
    assign out318 = tmp[318][STEP][0];
    assign out319 = tmp[319][STEP][0];
    assign out320 = tmp[320][STEP][0];
    assign out321 = tmp[321][STEP][0];
    assign out322 = tmp[322][STEP][0];
    assign out323 = tmp[323][STEP][0];
    assign out324 = tmp[324][STEP][0];
    assign out325 = tmp[325][STEP][0];
    assign out326 = tmp[326][STEP][0];
    assign out327 = tmp[327][STEP][0];
    assign out328 = tmp[328][STEP][0];
    assign out329 = tmp[329][STEP][0];
    assign out330 = tmp[330][STEP][0];
    assign out331 = tmp[331][STEP][0];
    assign out332 = tmp[332][STEP][0];
    assign out333 = tmp[333][STEP][0];
    assign out334 = tmp[334][STEP][0];
    assign out335 = tmp[335][STEP][0];
    assign out336 = tmp[336][STEP][0];
    assign out337 = tmp[337][STEP][0];
    assign out338 = tmp[338][STEP][0];
    assign out339 = tmp[339][STEP][0];
    assign out340 = tmp[340][STEP][0];
    assign out341 = tmp[341][STEP][0];
    assign out342 = tmp[342][STEP][0];
    assign out343 = tmp[343][STEP][0];
    assign out344 = tmp[344][STEP][0];
    assign out345 = tmp[345][STEP][0];
    assign out346 = tmp[346][STEP][0];
    assign out347 = tmp[347][STEP][0];
    assign out348 = tmp[348][STEP][0];
    assign out349 = tmp[349][STEP][0];
    assign out350 = tmp[350][STEP][0];
    assign out351 = tmp[351][STEP][0];
    assign out352 = tmp[352][STEP][0];
    assign out353 = tmp[353][STEP][0];
    assign out354 = tmp[354][STEP][0];
    assign out355 = tmp[355][STEP][0];
    assign out356 = tmp[356][STEP][0];
    assign out357 = tmp[357][STEP][0];
    assign out358 = tmp[358][STEP][0];
    assign out359 = tmp[359][STEP][0];
    assign out360 = tmp[360][STEP][0];
    assign out361 = tmp[361][STEP][0];
    assign out362 = tmp[362][STEP][0];
    assign out363 = tmp[363][STEP][0];
    assign out364 = tmp[364][STEP][0];
    assign out365 = tmp[365][STEP][0];
    assign out366 = tmp[366][STEP][0];
    assign out367 = tmp[367][STEP][0];
    assign out368 = tmp[368][STEP][0];
    assign out369 = tmp[369][STEP][0];
    assign out370 = tmp[370][STEP][0];
    assign out371 = tmp[371][STEP][0];
    assign out372 = tmp[372][STEP][0];
    assign out373 = tmp[373][STEP][0];
    assign out374 = tmp[374][STEP][0];
    assign out375 = tmp[375][STEP][0];
    assign out376 = tmp[376][STEP][0];
    assign out377 = tmp[377][STEP][0];
    assign out378 = tmp[378][STEP][0];
    assign out379 = tmp[379][STEP][0];
    assign out380 = tmp[380][STEP][0];
    assign out381 = tmp[381][STEP][0];
    assign out382 = tmp[382][STEP][0];
    assign out383 = tmp[383][STEP][0];
    assign out384 = tmp[384][STEP][0];
    assign out385 = tmp[385][STEP][0];
    assign out386 = tmp[386][STEP][0];
    assign out387 = tmp[387][STEP][0];
    assign out388 = tmp[388][STEP][0];
    assign out389 = tmp[389][STEP][0];
    assign out390 = tmp[390][STEP][0];
    assign out391 = tmp[391][STEP][0];
    assign out392 = tmp[392][STEP][0];
    assign out393 = tmp[393][STEP][0];
    assign out394 = tmp[394][STEP][0];
    assign out395 = tmp[395][STEP][0];
    assign out396 = tmp[396][STEP][0];
    assign out397 = tmp[397][STEP][0];
    assign out398 = tmp[398][STEP][0];
    assign out399 = tmp[399][STEP][0];
    assign out400 = tmp[400][STEP][0];
    assign out401 = tmp[401][STEP][0];
    assign out402 = tmp[402][STEP][0];
    assign out403 = tmp[403][STEP][0];
    assign out404 = tmp[404][STEP][0];
    assign out405 = tmp[405][STEP][0];
    assign out406 = tmp[406][STEP][0];
    assign out407 = tmp[407][STEP][0];
    assign out408 = tmp[408][STEP][0];
    assign out409 = tmp[409][STEP][0];
    assign out410 = tmp[410][STEP][0];
    assign out411 = tmp[411][STEP][0];
    assign out412 = tmp[412][STEP][0];
    assign out413 = tmp[413][STEP][0];
    assign out414 = tmp[414][STEP][0];
    assign out415 = tmp[415][STEP][0];
    assign out416 = tmp[416][STEP][0];
    assign out417 = tmp[417][STEP][0];
    assign out418 = tmp[418][STEP][0];
    assign out419 = tmp[419][STEP][0];
    assign out420 = tmp[420][STEP][0];
    assign out421 = tmp[421][STEP][0];
    assign out422 = tmp[422][STEP][0];
    assign out423 = tmp[423][STEP][0];
    assign out424 = tmp[424][STEP][0];
    assign out425 = tmp[425][STEP][0];
    assign out426 = tmp[426][STEP][0];
    assign out427 = tmp[427][STEP][0];
    assign out428 = tmp[428][STEP][0];
    assign out429 = tmp[429][STEP][0];
    assign out430 = tmp[430][STEP][0];
    assign out431 = tmp[431][STEP][0];
    assign out432 = tmp[432][STEP][0];
    assign out433 = tmp[433][STEP][0];
    assign out434 = tmp[434][STEP][0];
    assign out435 = tmp[435][STEP][0];
    assign out436 = tmp[436][STEP][0];
    assign out437 = tmp[437][STEP][0];
    assign out438 = tmp[438][STEP][0];
    assign out439 = tmp[439][STEP][0];
    assign out440 = tmp[440][STEP][0];
    assign out441 = tmp[441][STEP][0];
    assign out442 = tmp[442][STEP][0];
    assign out443 = tmp[443][STEP][0];
    assign out444 = tmp[444][STEP][0];
    assign out445 = tmp[445][STEP][0];
    assign out446 = tmp[446][STEP][0];
    assign out447 = tmp[447][STEP][0];
    assign out448 = tmp[448][STEP][0];
    assign out449 = tmp[449][STEP][0];
    assign out450 = tmp[450][STEP][0];
    assign out451 = tmp[451][STEP][0];
    assign out452 = tmp[452][STEP][0];
    assign out453 = tmp[453][STEP][0];
    assign out454 = tmp[454][STEP][0];
    assign out455 = tmp[455][STEP][0];
    assign out456 = tmp[456][STEP][0];
    assign out457 = tmp[457][STEP][0];
    assign out458 = tmp[458][STEP][0];
    assign out459 = tmp[459][STEP][0];
    assign out460 = tmp[460][STEP][0];
    assign out461 = tmp[461][STEP][0];
    assign out462 = tmp[462][STEP][0];
    assign out463 = tmp[463][STEP][0];
    assign out464 = tmp[464][STEP][0];
    assign out465 = tmp[465][STEP][0];
    assign out466 = tmp[466][STEP][0];
    assign out467 = tmp[467][STEP][0];
    assign out468 = tmp[468][STEP][0];
    assign out469 = tmp[469][STEP][0];
    assign out470 = tmp[470][STEP][0];
    assign out471 = tmp[471][STEP][0];
    assign out472 = tmp[472][STEP][0];
    assign out473 = tmp[473][STEP][0];
    assign out474 = tmp[474][STEP][0];
    assign out475 = tmp[475][STEP][0];
    assign out476 = tmp[476][STEP][0];
    assign out477 = tmp[477][STEP][0];
    assign out478 = tmp[478][STEP][0];
    assign out479 = tmp[479][STEP][0];
    assign out480 = tmp[480][STEP][0];
    assign out481 = tmp[481][STEP][0];
    assign out482 = tmp[482][STEP][0];
    assign out483 = tmp[483][STEP][0];
    assign out484 = tmp[484][STEP][0];
    assign out485 = tmp[485][STEP][0];
    assign out486 = tmp[486][STEP][0];
    assign out487 = tmp[487][STEP][0];
    assign out488 = tmp[488][STEP][0];
    assign out489 = tmp[489][STEP][0];
    assign out490 = tmp[490][STEP][0];
    assign out491 = tmp[491][STEP][0];
    assign out492 = tmp[492][STEP][0];
    assign out493 = tmp[493][STEP][0];
    assign out494 = tmp[494][STEP][0];
    assign out495 = tmp[495][STEP][0];
    assign out496 = tmp[496][STEP][0];
    assign out497 = tmp[497][STEP][0];
    assign out498 = tmp[498][STEP][0];
    assign out499 = tmp[499][STEP][0];
    assign out500 = tmp[500][STEP][0];
    assign out501 = tmp[501][STEP][0];
    assign out502 = tmp[502][STEP][0];
    assign out503 = tmp[503][STEP][0];
    assign out504 = tmp[504][STEP][0];
    assign out505 = tmp[505][STEP][0];
    assign out506 = tmp[506][STEP][0];
    assign out507 = tmp[507][STEP][0];
    assign out508 = tmp[508][STEP][0];
    assign out509 = tmp[509][STEP][0];
    assign out510 = tmp[510][STEP][0];
    assign out511 = tmp[511][STEP][0];
    assign out512 = tmp[512][STEP][0];
    assign out513 = tmp[513][STEP][0];
    assign out514 = tmp[514][STEP][0];
    assign out515 = tmp[515][STEP][0];
    assign out516 = tmp[516][STEP][0];
    assign out517 = tmp[517][STEP][0];
    assign out518 = tmp[518][STEP][0];
    assign out519 = tmp[519][STEP][0];
    assign out520 = tmp[520][STEP][0];
    assign out521 = tmp[521][STEP][0];
    assign out522 = tmp[522][STEP][0];
    assign out523 = tmp[523][STEP][0];
    assign out524 = tmp[524][STEP][0];
    assign out525 = tmp[525][STEP][0];
    assign out526 = tmp[526][STEP][0];
    assign out527 = tmp[527][STEP][0];
    assign out528 = tmp[528][STEP][0];
    assign out529 = tmp[529][STEP][0];
    assign out530 = tmp[530][STEP][0];
    assign out531 = tmp[531][STEP][0];
    assign out532 = tmp[532][STEP][0];
    assign out533 = tmp[533][STEP][0];
    assign out534 = tmp[534][STEP][0];
    assign out535 = tmp[535][STEP][0];
    assign out536 = tmp[536][STEP][0];
    assign out537 = tmp[537][STEP][0];
    assign out538 = tmp[538][STEP][0];
    assign out539 = tmp[539][STEP][0];
    assign out540 = tmp[540][STEP][0];
    assign out541 = tmp[541][STEP][0];
    assign out542 = tmp[542][STEP][0];
    assign out543 = tmp[543][STEP][0];
    assign out544 = tmp[544][STEP][0];
    assign out545 = tmp[545][STEP][0];
    assign out546 = tmp[546][STEP][0];
    assign out547 = tmp[547][STEP][0];
    assign out548 = tmp[548][STEP][0];
    assign out549 = tmp[549][STEP][0];
    assign out550 = tmp[550][STEP][0];
    assign out551 = tmp[551][STEP][0];
    assign out552 = tmp[552][STEP][0];
    assign out553 = tmp[553][STEP][0];
    assign out554 = tmp[554][STEP][0];
    assign out555 = tmp[555][STEP][0];
    assign out556 = tmp[556][STEP][0];
    assign out557 = tmp[557][STEP][0];
    assign out558 = tmp[558][STEP][0];
    assign out559 = tmp[559][STEP][0];
    assign out560 = tmp[560][STEP][0];
    assign out561 = tmp[561][STEP][0];
    assign out562 = tmp[562][STEP][0];
    assign out563 = tmp[563][STEP][0];
    assign out564 = tmp[564][STEP][0];
    assign out565 = tmp[565][STEP][0];
    assign out566 = tmp[566][STEP][0];
    assign out567 = tmp[567][STEP][0];
    assign out568 = tmp[568][STEP][0];
    assign out569 = tmp[569][STEP][0];
    assign out570 = tmp[570][STEP][0];
    assign out571 = tmp[571][STEP][0];
    assign out572 = tmp[572][STEP][0];
    assign out573 = tmp[573][STEP][0];
    assign out574 = tmp[574][STEP][0];
    assign out575 = tmp[575][STEP][0];
    assign out576 = tmp[576][STEP][0];
    assign out577 = tmp[577][STEP][0];
    assign out578 = tmp[578][STEP][0];
    assign out579 = tmp[579][STEP][0];
    assign out580 = tmp[580][STEP][0];
    assign out581 = tmp[581][STEP][0];
    assign out582 = tmp[582][STEP][0];
    assign out583 = tmp[583][STEP][0];
    assign out584 = tmp[584][STEP][0];
    assign out585 = tmp[585][STEP][0];
    assign out586 = tmp[586][STEP][0];
    assign out587 = tmp[587][STEP][0];
    assign out588 = tmp[588][STEP][0];
    assign out589 = tmp[589][STEP][0];
    assign out590 = tmp[590][STEP][0];
    assign out591 = tmp[591][STEP][0];
    assign out592 = tmp[592][STEP][0];
    assign out593 = tmp[593][STEP][0];
    assign out594 = tmp[594][STEP][0];
    assign out595 = tmp[595][STEP][0];
    assign out596 = tmp[596][STEP][0];
    assign out597 = tmp[597][STEP][0];
    assign out598 = tmp[598][STEP][0];
    assign out599 = tmp[599][STEP][0];
    assign out600 = tmp[600][STEP][0];
    assign out601 = tmp[601][STEP][0];
    assign out602 = tmp[602][STEP][0];
    assign out603 = tmp[603][STEP][0];
    assign out604 = tmp[604][STEP][0];
    assign out605 = tmp[605][STEP][0];
    assign out606 = tmp[606][STEP][0];
    assign out607 = tmp[607][STEP][0];
    assign out608 = tmp[608][STEP][0];
    assign out609 = tmp[609][STEP][0];
    assign out610 = tmp[610][STEP][0];
    assign out611 = tmp[611][STEP][0];
    assign out612 = tmp[612][STEP][0];
    assign out613 = tmp[613][STEP][0];
    assign out614 = tmp[614][STEP][0];
    assign out615 = tmp[615][STEP][0];
    assign out616 = tmp[616][STEP][0];
    assign out617 = tmp[617][STEP][0];
    assign out618 = tmp[618][STEP][0];
    assign out619 = tmp[619][STEP][0];
    assign out620 = tmp[620][STEP][0];
    assign out621 = tmp[621][STEP][0];
    assign out622 = tmp[622][STEP][0];
    assign out623 = tmp[623][STEP][0];
    assign out624 = tmp[624][STEP][0];
    assign out625 = tmp[625][STEP][0];
    assign out626 = tmp[626][STEP][0];
    assign out627 = tmp[627][STEP][0];
    assign out628 = tmp[628][STEP][0];
    assign out629 = tmp[629][STEP][0];
    assign out630 = tmp[630][STEP][0];
    assign out631 = tmp[631][STEP][0];
    assign out632 = tmp[632][STEP][0];
    assign out633 = tmp[633][STEP][0];
    assign out634 = tmp[634][STEP][0];
    assign out635 = tmp[635][STEP][0];
    assign out636 = tmp[636][STEP][0];
    assign out637 = tmp[637][STEP][0];
    assign out638 = tmp[638][STEP][0];
    assign out639 = tmp[639][STEP][0];
    assign out640 = tmp[640][STEP][0];
    assign out641 = tmp[641][STEP][0];
    assign out642 = tmp[642][STEP][0];
    assign out643 = tmp[643][STEP][0];
    assign out644 = tmp[644][STEP][0];
    assign out645 = tmp[645][STEP][0];
    assign out646 = tmp[646][STEP][0];
    assign out647 = tmp[647][STEP][0];
    assign out648 = tmp[648][STEP][0];
    assign out649 = tmp[649][STEP][0];
    assign out650 = tmp[650][STEP][0];
    assign out651 = tmp[651][STEP][0];
    assign out652 = tmp[652][STEP][0];
    assign out653 = tmp[653][STEP][0];
    assign out654 = tmp[654][STEP][0];
    assign out655 = tmp[655][STEP][0];
    assign out656 = tmp[656][STEP][0];
    assign out657 = tmp[657][STEP][0];
    assign out658 = tmp[658][STEP][0];
    assign out659 = tmp[659][STEP][0];
    assign out660 = tmp[660][STEP][0];
    assign out661 = tmp[661][STEP][0];
    assign out662 = tmp[662][STEP][0];
    assign out663 = tmp[663][STEP][0];
    assign out664 = tmp[664][STEP][0];
    assign out665 = tmp[665][STEP][0];
    assign out666 = tmp[666][STEP][0];
    assign out667 = tmp[667][STEP][0];
    assign out668 = tmp[668][STEP][0];
    assign out669 = tmp[669][STEP][0];
    assign out670 = tmp[670][STEP][0];
    assign out671 = tmp[671][STEP][0];
    assign out672 = tmp[672][STEP][0];
    assign out673 = tmp[673][STEP][0];
    assign out674 = tmp[674][STEP][0];
    assign out675 = tmp[675][STEP][0];
    assign out676 = tmp[676][STEP][0];
    assign out677 = tmp[677][STEP][0];
    assign out678 = tmp[678][STEP][0];
    assign out679 = tmp[679][STEP][0];
    assign out680 = tmp[680][STEP][0];
    assign out681 = tmp[681][STEP][0];
    assign out682 = tmp[682][STEP][0];
    assign out683 = tmp[683][STEP][0];
    assign out684 = tmp[684][STEP][0];
    assign out685 = tmp[685][STEP][0];
    assign out686 = tmp[686][STEP][0];
    assign out687 = tmp[687][STEP][0];
    assign out688 = tmp[688][STEP][0];
    assign out689 = tmp[689][STEP][0];
    assign out690 = tmp[690][STEP][0];
    assign out691 = tmp[691][STEP][0];
    assign out692 = tmp[692][STEP][0];
    assign out693 = tmp[693][STEP][0];
    assign out694 = tmp[694][STEP][0];
    assign out695 = tmp[695][STEP][0];
    assign out696 = tmp[696][STEP][0];
    assign out697 = tmp[697][STEP][0];
    assign out698 = tmp[698][STEP][0];
    assign out699 = tmp[699][STEP][0];
    assign out700 = tmp[700][STEP][0];
    assign out701 = tmp[701][STEP][0];
    assign out702 = tmp[702][STEP][0];
    assign out703 = tmp[703][STEP][0];
    assign out704 = tmp[704][STEP][0];
    assign out705 = tmp[705][STEP][0];
    assign out706 = tmp[706][STEP][0];
    assign out707 = tmp[707][STEP][0];
    assign out708 = tmp[708][STEP][0];
    assign out709 = tmp[709][STEP][0];
    assign out710 = tmp[710][STEP][0];
    assign out711 = tmp[711][STEP][0];
    assign out712 = tmp[712][STEP][0];
    assign out713 = tmp[713][STEP][0];
    assign out714 = tmp[714][STEP][0];
    assign out715 = tmp[715][STEP][0];
    assign out716 = tmp[716][STEP][0];
    assign out717 = tmp[717][STEP][0];
    assign out718 = tmp[718][STEP][0];
    assign out719 = tmp[719][STEP][0];
    assign out720 = tmp[720][STEP][0];
    assign out721 = tmp[721][STEP][0];
    assign out722 = tmp[722][STEP][0];
    assign out723 = tmp[723][STEP][0];
    assign out724 = tmp[724][STEP][0];
    assign out725 = tmp[725][STEP][0];
    assign out726 = tmp[726][STEP][0];
    assign out727 = tmp[727][STEP][0];
    assign out728 = tmp[728][STEP][0];
    assign out729 = tmp[729][STEP][0];
    assign out730 = tmp[730][STEP][0];
    assign out731 = tmp[731][STEP][0];
    assign out732 = tmp[732][STEP][0];
    assign out733 = tmp[733][STEP][0];
    assign out734 = tmp[734][STEP][0];
    assign out735 = tmp[735][STEP][0];
    assign out736 = tmp[736][STEP][0];
    assign out737 = tmp[737][STEP][0];
    assign out738 = tmp[738][STEP][0];
    assign out739 = tmp[739][STEP][0];
    assign out740 = tmp[740][STEP][0];
    assign out741 = tmp[741][STEP][0];
    assign out742 = tmp[742][STEP][0];
    assign out743 = tmp[743][STEP][0];
    assign out744 = tmp[744][STEP][0];
    assign out745 = tmp[745][STEP][0];
    assign out746 = tmp[746][STEP][0];
    assign out747 = tmp[747][STEP][0];
    assign out748 = tmp[748][STEP][0];
    assign out749 = tmp[749][STEP][0];
    assign out750 = tmp[750][STEP][0];
    assign out751 = tmp[751][STEP][0];
    assign out752 = tmp[752][STEP][0];
    assign out753 = tmp[753][STEP][0];
    assign out754 = tmp[754][STEP][0];
    assign out755 = tmp[755][STEP][0];
    assign out756 = tmp[756][STEP][0];
    assign out757 = tmp[757][STEP][0];
    assign out758 = tmp[758][STEP][0];
    assign out759 = tmp[759][STEP][0];
    assign out760 = tmp[760][STEP][0];
    assign out761 = tmp[761][STEP][0];
    assign out762 = tmp[762][STEP][0];
    assign out763 = tmp[763][STEP][0];
    assign out764 = tmp[764][STEP][0];
    assign out765 = tmp[765][STEP][0];
    assign out766 = tmp[766][STEP][0];
    assign out767 = tmp[767][STEP][0];
    assign out768 = tmp[768][STEP][0];
    assign out769 = tmp[769][STEP][0];
    assign out770 = tmp[770][STEP][0];
    assign out771 = tmp[771][STEP][0];
    assign out772 = tmp[772][STEP][0];
    assign out773 = tmp[773][STEP][0];
    assign out774 = tmp[774][STEP][0];
    assign out775 = tmp[775][STEP][0];
    assign out776 = tmp[776][STEP][0];
    assign out777 = tmp[777][STEP][0];
    assign out778 = tmp[778][STEP][0];
    assign out779 = tmp[779][STEP][0];
    assign out780 = tmp[780][STEP][0];
    assign out781 = tmp[781][STEP][0];
    assign out782 = tmp[782][STEP][0];
    assign out783 = tmp[783][STEP][0];
    assign out784 = tmp[784][STEP][0];
    assign out785 = tmp[785][STEP][0];
    assign out786 = tmp[786][STEP][0];
    assign out787 = tmp[787][STEP][0];
    assign out788 = tmp[788][STEP][0];
    assign out789 = tmp[789][STEP][0];
    assign out790 = tmp[790][STEP][0];
    assign out791 = tmp[791][STEP][0];
    assign out792 = tmp[792][STEP][0];
    assign out793 = tmp[793][STEP][0];
    assign out794 = tmp[794][STEP][0];
    assign out795 = tmp[795][STEP][0];
    assign out796 = tmp[796][STEP][0];
    assign out797 = tmp[797][STEP][0];
    assign out798 = tmp[798][STEP][0];
    assign out799 = tmp[799][STEP][0];
    assign out800 = tmp[800][STEP][0];
    assign out801 = tmp[801][STEP][0];
    assign out802 = tmp[802][STEP][0];
    assign out803 = tmp[803][STEP][0];
    assign out804 = tmp[804][STEP][0];
    assign out805 = tmp[805][STEP][0];
    assign out806 = tmp[806][STEP][0];
    assign out807 = tmp[807][STEP][0];
    assign out808 = tmp[808][STEP][0];
    assign out809 = tmp[809][STEP][0];
    assign out810 = tmp[810][STEP][0];
    assign out811 = tmp[811][STEP][0];
    assign out812 = tmp[812][STEP][0];
    assign out813 = tmp[813][STEP][0];
    assign out814 = tmp[814][STEP][0];
    assign out815 = tmp[815][STEP][0];
    assign out816 = tmp[816][STEP][0];
    assign out817 = tmp[817][STEP][0];
    assign out818 = tmp[818][STEP][0];
    assign out819 = tmp[819][STEP][0];
    assign out820 = tmp[820][STEP][0];
    assign out821 = tmp[821][STEP][0];
    assign out822 = tmp[822][STEP][0];
    assign out823 = tmp[823][STEP][0];
    assign out824 = tmp[824][STEP][0];
    assign out825 = tmp[825][STEP][0];
    assign out826 = tmp[826][STEP][0];
    assign out827 = tmp[827][STEP][0];
    assign out828 = tmp[828][STEP][0];
    assign out829 = tmp[829][STEP][0];
    assign out830 = tmp[830][STEP][0];
    assign out831 = tmp[831][STEP][0];
    assign out832 = tmp[832][STEP][0];
    assign out833 = tmp[833][STEP][0];
    assign out834 = tmp[834][STEP][0];
    assign out835 = tmp[835][STEP][0];
    assign out836 = tmp[836][STEP][0];
    assign out837 = tmp[837][STEP][0];
    assign out838 = tmp[838][STEP][0];
    assign out839 = tmp[839][STEP][0];
    assign out840 = tmp[840][STEP][0];
    assign out841 = tmp[841][STEP][0];
    assign out842 = tmp[842][STEP][0];
    assign out843 = tmp[843][STEP][0];
    assign out844 = tmp[844][STEP][0];
    assign out845 = tmp[845][STEP][0];
    assign out846 = tmp[846][STEP][0];
    assign out847 = tmp[847][STEP][0];
    assign out848 = tmp[848][STEP][0];
    assign out849 = tmp[849][STEP][0];
    assign out850 = tmp[850][STEP][0];
    assign out851 = tmp[851][STEP][0];
    assign out852 = tmp[852][STEP][0];
    assign out853 = tmp[853][STEP][0];
    assign out854 = tmp[854][STEP][0];
    assign out855 = tmp[855][STEP][0];
    assign out856 = tmp[856][STEP][0];
    assign out857 = tmp[857][STEP][0];
    assign out858 = tmp[858][STEP][0];
    assign out859 = tmp[859][STEP][0];
    assign out860 = tmp[860][STEP][0];
    assign out861 = tmp[861][STEP][0];
    assign out862 = tmp[862][STEP][0];
    assign out863 = tmp[863][STEP][0];
    assign out864 = tmp[864][STEP][0];
    assign out865 = tmp[865][STEP][0];
    assign out866 = tmp[866][STEP][0];
    assign out867 = tmp[867][STEP][0];
    assign out868 = tmp[868][STEP][0];
    assign out869 = tmp[869][STEP][0];
    assign out870 = tmp[870][STEP][0];
    assign out871 = tmp[871][STEP][0];
    assign out872 = tmp[872][STEP][0];
    assign out873 = tmp[873][STEP][0];
    assign out874 = tmp[874][STEP][0];
    assign out875 = tmp[875][STEP][0];
    assign out876 = tmp[876][STEP][0];
    assign out877 = tmp[877][STEP][0];
    assign out878 = tmp[878][STEP][0];
    assign out879 = tmp[879][STEP][0];
    assign out880 = tmp[880][STEP][0];
    assign out881 = tmp[881][STEP][0];
    assign out882 = tmp[882][STEP][0];
    assign out883 = tmp[883][STEP][0];
    assign out884 = tmp[884][STEP][0];
    assign out885 = tmp[885][STEP][0];
    assign out886 = tmp[886][STEP][0];
    assign out887 = tmp[887][STEP][0];
    assign out888 = tmp[888][STEP][0];
    assign out889 = tmp[889][STEP][0];
    assign out890 = tmp[890][STEP][0];
    assign out891 = tmp[891][STEP][0];
    assign out892 = tmp[892][STEP][0];
    assign out893 = tmp[893][STEP][0];
    assign out894 = tmp[894][STEP][0];
    assign out895 = tmp[895][STEP][0];
    assign out896 = tmp[896][STEP][0];
    assign out897 = tmp[897][STEP][0];
    assign out898 = tmp[898][STEP][0];
    assign out899 = tmp[899][STEP][0];
    assign out900 = tmp[900][STEP][0];
    assign out901 = tmp[901][STEP][0];
    assign out902 = tmp[902][STEP][0];
    assign out903 = tmp[903][STEP][0];
    assign out904 = tmp[904][STEP][0];
    assign out905 = tmp[905][STEP][0];
    assign out906 = tmp[906][STEP][0];
    assign out907 = tmp[907][STEP][0];
    assign out908 = tmp[908][STEP][0];
    assign out909 = tmp[909][STEP][0];
    assign out910 = tmp[910][STEP][0];
    assign out911 = tmp[911][STEP][0];
    assign out912 = tmp[912][STEP][0];
    assign out913 = tmp[913][STEP][0];
    assign out914 = tmp[914][STEP][0];
    assign out915 = tmp[915][STEP][0];
    assign out916 = tmp[916][STEP][0];
    assign out917 = tmp[917][STEP][0];
    assign out918 = tmp[918][STEP][0];
    assign out919 = tmp[919][STEP][0];
    assign out920 = tmp[920][STEP][0];
    assign out921 = tmp[921][STEP][0];
    assign out922 = tmp[922][STEP][0];
    assign out923 = tmp[923][STEP][0];
    assign out924 = tmp[924][STEP][0];
    assign out925 = tmp[925][STEP][0];
    assign out926 = tmp[926][STEP][0];
    assign out927 = tmp[927][STEP][0];
    assign out928 = tmp[928][STEP][0];
    assign out929 = tmp[929][STEP][0];
    assign out930 = tmp[930][STEP][0];
    assign out931 = tmp[931][STEP][0];
    assign out932 = tmp[932][STEP][0];
    assign out933 = tmp[933][STEP][0];
    assign out934 = tmp[934][STEP][0];
    assign out935 = tmp[935][STEP][0];
    assign out936 = tmp[936][STEP][0];
    assign out937 = tmp[937][STEP][0];
    assign out938 = tmp[938][STEP][0];
    assign out939 = tmp[939][STEP][0];
    assign out940 = tmp[940][STEP][0];
    assign out941 = tmp[941][STEP][0];
    assign out942 = tmp[942][STEP][0];
    assign out943 = tmp[943][STEP][0];
    assign out944 = tmp[944][STEP][0];
    assign out945 = tmp[945][STEP][0];
    assign out946 = tmp[946][STEP][0];
    assign out947 = tmp[947][STEP][0];
    assign out948 = tmp[948][STEP][0];
    assign out949 = tmp[949][STEP][0];
    assign out950 = tmp[950][STEP][0];
    assign out951 = tmp[951][STEP][0];
    assign out952 = tmp[952][STEP][0];
    assign out953 = tmp[953][STEP][0];
    assign out954 = tmp[954][STEP][0];
    assign out955 = tmp[955][STEP][0];
    assign out956 = tmp[956][STEP][0];
    assign out957 = tmp[957][STEP][0];
    assign out958 = tmp[958][STEP][0];
    assign out959 = tmp[959][STEP][0];
    assign out960 = tmp[960][STEP][0];
    assign out961 = tmp[961][STEP][0];
    assign out962 = tmp[962][STEP][0];
    assign out963 = tmp[963][STEP][0];
    assign out964 = tmp[964][STEP][0];
    assign out965 = tmp[965][STEP][0];
    assign out966 = tmp[966][STEP][0];
    assign out967 = tmp[967][STEP][0];
    assign out968 = tmp[968][STEP][0];
    assign out969 = tmp[969][STEP][0];
    assign out970 = tmp[970][STEP][0];
    assign out971 = tmp[971][STEP][0];
    assign out972 = tmp[972][STEP][0];
    assign out973 = tmp[973][STEP][0];
    assign out974 = tmp[974][STEP][0];
    assign out975 = tmp[975][STEP][0];
    assign out976 = tmp[976][STEP][0];
    assign out977 = tmp[977][STEP][0];
    assign out978 = tmp[978][STEP][0];
    assign out979 = tmp[979][STEP][0];
    assign out980 = tmp[980][STEP][0];
    assign out981 = tmp[981][STEP][0];
    assign out982 = tmp[982][STEP][0];
    assign out983 = tmp[983][STEP][0];
    assign out984 = tmp[984][STEP][0];
    assign out985 = tmp[985][STEP][0];
    assign out986 = tmp[986][STEP][0];
    assign out987 = tmp[987][STEP][0];
    assign out988 = tmp[988][STEP][0];
    assign out989 = tmp[989][STEP][0];
    assign out990 = tmp[990][STEP][0];
    assign out991 = tmp[991][STEP][0];
    assign out992 = tmp[992][STEP][0];
    assign out993 = tmp[993][STEP][0];
    assign out994 = tmp[994][STEP][0];
    assign out995 = tmp[995][STEP][0];
    assign out996 = tmp[996][STEP][0];
    assign out997 = tmp[997][STEP][0];
    assign out998 = tmp[998][STEP][0];
    assign out999 = tmp[999][STEP][0];
    assign out1000 = tmp[1000][STEP][0];
    assign out1001 = tmp[1001][STEP][0];
    assign out1002 = tmp[1002][STEP][0];
    assign out1003 = tmp[1003][STEP][0];
    assign out1004 = tmp[1004][STEP][0];
    assign out1005 = tmp[1005][STEP][0];
    assign out1006 = tmp[1006][STEP][0];
    assign out1007 = tmp[1007][STEP][0];
    assign out1008 = tmp[1008][STEP][0];
    assign out1009 = tmp[1009][STEP][0];
    assign out1010 = tmp[1010][STEP][0];
    assign out1011 = tmp[1011][STEP][0];
    assign out1012 = tmp[1012][STEP][0];
    assign out1013 = tmp[1013][STEP][0];
    assign out1014 = tmp[1014][STEP][0];
    assign out1015 = tmp[1015][STEP][0];
    assign out1016 = tmp[1016][STEP][0];
    assign out1017 = tmp[1017][STEP][0];
    assign out1018 = tmp[1018][STEP][0];
    assign out1019 = tmp[1019][STEP][0];
    assign out1020 = tmp[1020][STEP][0];
    assign out1021 = tmp[1021][STEP][0];
    assign out1022 = tmp[1022][STEP][0];
    assign out1023 = tmp[1023][STEP][0];
        /*
    initial begin
        #20000
        
        for (y = 0; y < STEP; y = y + 1)begin
            for (x = 0; x < N/2; x=x+1)begin
                $display("tmp[%d*2][%d][0]=%x\n",x,y,tmp[x*2][y][0]);
                $display("tmp[%d+4][2-%d][1]=%x\n",x,y,tmp[x+4][2-y][1]);
                $display("tmp[%d*2+1][%d][0]=%x\n",x,y,tmp[x*2+1][y][0]);
                $display("w[%d][%d][0]=%x\n\n",x,y,w[x][y][0]);
                $display("tmp[%d][%d+1][0]=%x\n\n",x,y,tmp[x][y+1][0]);
            end
            for (x = 0; x < N/2; x=x+1)begin
                $display("tmp[%d][2-%d][1]=%x\n",x,y,tmp[x][2-y][1]);
                $display("tmp[%d*2][%d][0]=%x\n",x,y,tmp[x*2][y][0]);
                $display("tmp[%d*2+1][%d][0]=%x\n",x,y,tmp[x*2+1][y][0]);
                $display("w[%d+4][%d][0]=%x\n\n",x,y,w[x+4][y][0]);
                $display("tmp[%d+4][%d+1][0]=%x\n\n",x,y,tmp[x+4][y+1][0]);
            end
        end
        for (y = 0; y < STEP; y = y + 1)begin
            $display("-------------------------------%d---------------",y);
            for (x = 0; x < N/2; x=x+1)begin
                $display("tmp[%d][%d][1]=%x\n",x,y,tmp[x][y][1]);
                $display("tmp[%d+4][%d][1]=%x\n",x,y,tmp[x+4][y][1]);
                $display("tmp[%d*2+1][2-%d][0]=%x\n",x,y,tmp[x*2+1][2-y][0]);
                $display("w[%d*2][%d][1]=%x\n\n",x,y,w[x*2][y][1]);
                #5
                $display("tmp[%d*2][%d+1][1]=%x\n\n",x,y,tmp[x*2][y+1][1]);
            end
            for (x = 0; x < N/2; x=x+1)begin
                $display("tmp[%d][%d][1]=%x\n",x,y,tmp[x][y][1]);
                $display("tmp[%d*2][2-%d][0]=%x\n",x,y,tmp[x*2][2-y][0]);
                $display("tmp[%d+4][%d][1]=%x\n",x,y,tmp[x+4][y][1]);
                $display("w[%d*2+1][%d][1]=%x\n\n",x,y,w[x*2+1][y][1]);
                #5
                $display("tmp[%d*2+1][%d+1][1]=%x\n\n",x,y,tmp[x*2+1][y+1][1]);
            end
        end
    end
        */

    generate
        for(j = 0; j < STEP; j = j +1)
            for(i = 0; i < N/2; i = i + 1)begin
                cal1 l1(tmp[i*2][j][0],tmp[i+N/2][STEP-1-j][1],tmp[i*2+1][j][0],w[i][j][0]);
                cal2 l2(tmp[i][STEP-1-j][1],tmp[i*2][j][0],tmp[i*2+1][j][0],w[i+N/2][j][0]);
            end
        for(j = 0; j < STEP; j = j +1)
            for(i = 0; i < N/2; i = i + 1)begin
                cal1 r1(tmp[i][j][1],tmp[i+N/2][j][1],tmp[i*2+1][STEP-1-j][0],w[i*2][j][1]);
                cal2 r2(tmp[i][j][1],tmp[i*2][STEP-1-j][0],tmp[i+N/2][j][1],w[i*2+1][j][1]);
            end
    endgenerate

    always@(posedge clk, negedge rst_n)begin
        if(!rst_n)begin
            stage <= 4'd0;
            done <= 1'd0;
            counter <= 4'd0;
            for (x = 0; x < N; x = x + 1)
                for (y = 1; y <= STEP; y = y + 1)
                    for (z = 0; z < 2; z = z + 1)
                        tmp[x][y][z] <= `_SIZE'd0;
            tmp[0][0][1] <= 20'h00000;
            tmp[1][0][1] <= 20'h00000;
            tmp[2][0][1] <= 20'h00000;
            tmp[3][0][1] <= 20'h00000;
            tmp[4][0][1] <= 20'h00000;
            tmp[5][0][1] <= 20'h00000;
            tmp[6][0][1] <= 20'h00000;
            tmp[7][0][1] <= 20'h00000;
            tmp[8][0][1] <= 20'h00000;
            tmp[9][0][1] <= 20'h00000;
            tmp[10][0][1] <= 20'h00000;
            tmp[11][0][1] <= 20'h00000;
            tmp[12][0][1] <= 20'h00000;
            tmp[13][0][1] <= 20'h00000;
            tmp[14][0][1] <= 20'h00000;
            tmp[15][0][1] <= 20'h7ffff;
            tmp[16][0][1] <= 20'h00000;
            tmp[17][0][1] <= 20'h00000;
            tmp[18][0][1] <= 20'h00000;
            tmp[19][0][1] <= 20'h00000;
            tmp[20][0][1] <= 20'h00000;
            tmp[21][0][1] <= 20'h00000;
            tmp[22][0][1] <= 20'h00000;
            tmp[23][0][1] <= 20'h7ffff;
            tmp[24][0][1] <= 20'h00000;
            tmp[25][0][1] <= 20'h00000;
            tmp[26][0][1] <= 20'h00000;
            tmp[27][0][1] <= 20'h7ffff;
            tmp[28][0][1] <= 20'h00000;
            tmp[29][0][1] <= 20'h00000;
            tmp[30][0][1] <= 20'h00000;
            tmp[31][0][1] <= 20'h7ffff;
            tmp[32][0][1] <= 20'h00000;
            tmp[33][0][1] <= 20'h00000;
            tmp[34][0][1] <= 20'h00000;
            tmp[35][0][1] <= 20'h00000;
            tmp[36][0][1] <= 20'h00000;
            tmp[37][0][1] <= 20'h00000;
            tmp[38][0][1] <= 20'h00000;
            tmp[39][0][1] <= 20'h7ffff;
            tmp[40][0][1] <= 20'h00000;
            tmp[41][0][1] <= 20'h00000;
            tmp[42][0][1] <= 20'h00000;
            tmp[43][0][1] <= 20'h7ffff;
            tmp[44][0][1] <= 20'h00000;
            tmp[45][0][1] <= 20'h00000;
            tmp[46][0][1] <= 20'h00000;
            tmp[47][0][1] <= 20'h7ffff;
            tmp[48][0][1] <= 20'h00000;
            tmp[49][0][1] <= 20'h00000;
            tmp[50][0][1] <= 20'h00000;
            tmp[51][0][1] <= 20'h7ffff;
            tmp[52][0][1] <= 20'h00000;
            tmp[53][0][1] <= 20'h00000;
            tmp[54][0][1] <= 20'h00000;
            tmp[55][0][1] <= 20'h7ffff;
            tmp[56][0][1] <= 20'h00000;
            tmp[57][0][1] <= 20'h00000;
            tmp[58][0][1] <= 20'h00000;
            tmp[59][0][1] <= 20'h7ffff;
            tmp[60][0][1] <= 20'h00000;
            tmp[61][0][1] <= 20'h7ffff;
            tmp[62][0][1] <= 20'h7ffff;
            tmp[63][0][1] <= 20'h7ffff;
            tmp[64][0][1] <= 20'h00000;
            tmp[65][0][1] <= 20'h00000;
            tmp[66][0][1] <= 20'h00000;
            tmp[67][0][1] <= 20'h00000;
            tmp[68][0][1] <= 20'h00000;
            tmp[69][0][1] <= 20'h00000;
            tmp[70][0][1] <= 20'h00000;
            tmp[71][0][1] <= 20'h7ffff;
            tmp[72][0][1] <= 20'h00000;
            tmp[73][0][1] <= 20'h00000;
            tmp[74][0][1] <= 20'h00000;
            tmp[75][0][1] <= 20'h7ffff;
            tmp[76][0][1] <= 20'h00000;
            tmp[77][0][1] <= 20'h00000;
            tmp[78][0][1] <= 20'h00000;
            tmp[79][0][1] <= 20'h7ffff;
            tmp[80][0][1] <= 20'h00000;
            tmp[81][0][1] <= 20'h00000;
            tmp[82][0][1] <= 20'h00000;
            tmp[83][0][1] <= 20'h00000;
            tmp[84][0][1] <= 20'h00000;
            tmp[85][0][1] <= 20'h00000;
            tmp[86][0][1] <= 20'h00000;
            tmp[87][0][1] <= 20'h7ffff;
            tmp[88][0][1] <= 20'h00000;
            tmp[89][0][1] <= 20'h00000;
            tmp[90][0][1] <= 20'h00000;
            tmp[91][0][1] <= 20'h7ffff;
            tmp[92][0][1] <= 20'h00000;
            tmp[93][0][1] <= 20'h7ffff;
            tmp[94][0][1] <= 20'h7ffff;
            tmp[95][0][1] <= 20'h7ffff;
            tmp[96][0][1] <= 20'h00000;
            tmp[97][0][1] <= 20'h00000;
            tmp[98][0][1] <= 20'h00000;
            tmp[99][0][1] <= 20'h00000;
            tmp[100][0][1] <= 20'h00000;
            tmp[101][0][1] <= 20'h00000;
            tmp[102][0][1] <= 20'h00000;
            tmp[103][0][1] <= 20'h7ffff;
            tmp[104][0][1] <= 20'h00000;
            tmp[105][0][1] <= 20'h00000;
            tmp[106][0][1] <= 20'h00000;
            tmp[107][0][1] <= 20'h7ffff;
            tmp[108][0][1] <= 20'h00000;
            tmp[109][0][1] <= 20'h7ffff;
            tmp[110][0][1] <= 20'h7ffff;
            tmp[111][0][1] <= 20'h7ffff;
            tmp[112][0][1] <= 20'h00000;
            tmp[113][0][1] <= 20'h00000;
            tmp[114][0][1] <= 20'h00000;
            tmp[115][0][1] <= 20'h7ffff;
            tmp[116][0][1] <= 20'h00000;
            tmp[117][0][1] <= 20'h7ffff;
            tmp[118][0][1] <= 20'h7ffff;
            tmp[119][0][1] <= 20'h7ffff;
            tmp[120][0][1] <= 20'h00000;
            tmp[121][0][1] <= 20'h7ffff;
            tmp[122][0][1] <= 20'h7ffff;
            tmp[123][0][1] <= 20'h7ffff;
            tmp[124][0][1] <= 20'h00000;
            tmp[125][0][1] <= 20'h7ffff;
            tmp[126][0][1] <= 20'h7ffff;
            tmp[127][0][1] <= 20'h7ffff;
            tmp[128][0][1] <= 20'h00000;
            tmp[129][0][1] <= 20'h00000;
            tmp[130][0][1] <= 20'h00000;
            tmp[131][0][1] <= 20'h00000;
            tmp[132][0][1] <= 20'h00000;
            tmp[133][0][1] <= 20'h00000;
            tmp[134][0][1] <= 20'h00000;
            tmp[135][0][1] <= 20'h7ffff;
            tmp[136][0][1] <= 20'h00000;
            tmp[137][0][1] <= 20'h00000;
            tmp[138][0][1] <= 20'h00000;
            tmp[139][0][1] <= 20'h7ffff;
            tmp[140][0][1] <= 20'h00000;
            tmp[141][0][1] <= 20'h00000;
            tmp[142][0][1] <= 20'h00000;
            tmp[143][0][1] <= 20'h7ffff;
            tmp[144][0][1] <= 20'h00000;
            tmp[145][0][1] <= 20'h00000;
            tmp[146][0][1] <= 20'h00000;
            tmp[147][0][1] <= 20'h00000;
            tmp[148][0][1] <= 20'h00000;
            tmp[149][0][1] <= 20'h00000;
            tmp[150][0][1] <= 20'h00000;
            tmp[151][0][1] <= 20'h7ffff;
            tmp[152][0][1] <= 20'h00000;
            tmp[153][0][1] <= 20'h00000;
            tmp[154][0][1] <= 20'h00000;
            tmp[155][0][1] <= 20'h7ffff;
            tmp[156][0][1] <= 20'h00000;
            tmp[157][0][1] <= 20'h7ffff;
            tmp[158][0][1] <= 20'h7ffff;
            tmp[159][0][1] <= 20'h7ffff;
            tmp[160][0][1] <= 20'h00000;
            tmp[161][0][1] <= 20'h00000;
            tmp[162][0][1] <= 20'h00000;
            tmp[163][0][1] <= 20'h00000;
            tmp[164][0][1] <= 20'h00000;
            tmp[165][0][1] <= 20'h00000;
            tmp[166][0][1] <= 20'h00000;
            tmp[167][0][1] <= 20'h7ffff;
            tmp[168][0][1] <= 20'h00000;
            tmp[169][0][1] <= 20'h00000;
            tmp[170][0][1] <= 20'h00000;
            tmp[171][0][1] <= 20'h7ffff;
            tmp[172][0][1] <= 20'h00000;
            tmp[173][0][1] <= 20'h7ffff;
            tmp[174][0][1] <= 20'h7ffff;
            tmp[175][0][1] <= 20'h7ffff;
            tmp[176][0][1] <= 20'h00000;
            tmp[177][0][1] <= 20'h00000;
            tmp[178][0][1] <= 20'h00000;
            tmp[179][0][1] <= 20'h7ffff;
            tmp[180][0][1] <= 20'h00000;
            tmp[181][0][1] <= 20'h7ffff;
            tmp[182][0][1] <= 20'h7ffff;
            tmp[183][0][1] <= 20'h7ffff;
            tmp[184][0][1] <= 20'h00000;
            tmp[185][0][1] <= 20'h7ffff;
            tmp[186][0][1] <= 20'h7ffff;
            tmp[187][0][1] <= 20'h7ffff;
            tmp[188][0][1] <= 20'h00000;
            tmp[189][0][1] <= 20'h7ffff;
            tmp[190][0][1] <= 20'h7ffff;
            tmp[191][0][1] <= 20'h7ffff;
            tmp[192][0][1] <= 20'h00000;
            tmp[193][0][1] <= 20'h00000;
            tmp[194][0][1] <= 20'h00000;
            tmp[195][0][1] <= 20'h00000;
            tmp[196][0][1] <= 20'h00000;
            tmp[197][0][1] <= 20'h00000;
            tmp[198][0][1] <= 20'h00000;
            tmp[199][0][1] <= 20'h7ffff;
            tmp[200][0][1] <= 20'h00000;
            tmp[201][0][1] <= 20'h00000;
            tmp[202][0][1] <= 20'h00000;
            tmp[203][0][1] <= 20'h7ffff;
            tmp[204][0][1] <= 20'h00000;
            tmp[205][0][1] <= 20'h7ffff;
            tmp[206][0][1] <= 20'h7ffff;
            tmp[207][0][1] <= 20'h7ffff;
            tmp[208][0][1] <= 20'h00000;
            tmp[209][0][1] <= 20'h00000;
            tmp[210][0][1] <= 20'h00000;
            tmp[211][0][1] <= 20'h7ffff;
            tmp[212][0][1] <= 20'h00000;
            tmp[213][0][1] <= 20'h7ffff;
            tmp[214][0][1] <= 20'h7ffff;
            tmp[215][0][1] <= 20'h7ffff;
            tmp[216][0][1] <= 20'h00000;
            tmp[217][0][1] <= 20'h7ffff;
            tmp[218][0][1] <= 20'h00000;
            tmp[219][0][1] <= 20'h7ffff;
            tmp[220][0][1] <= 20'h00000;
            tmp[221][0][1] <= 20'h7ffff;
            tmp[222][0][1] <= 20'h7ffff;
            tmp[223][0][1] <= 20'h7ffff;
            tmp[224][0][1] <= 20'h00000;
            tmp[225][0][1] <= 20'h00000;
            tmp[226][0][1] <= 20'h00000;
            tmp[227][0][1] <= 20'h7ffff;
            tmp[228][0][1] <= 20'h00000;
            tmp[229][0][1] <= 20'h7ffff;
            tmp[230][0][1] <= 20'h7ffff;
            tmp[231][0][1] <= 20'h7ffff;
            tmp[232][0][1] <= 20'h00000;
            tmp[233][0][1] <= 20'h7ffff;
            tmp[234][0][1] <= 20'h00000;
            tmp[235][0][1] <= 20'h7ffff;
            tmp[236][0][1] <= 20'h00000;
            tmp[237][0][1] <= 20'h7ffff;
            tmp[238][0][1] <= 20'h7ffff;
            tmp[239][0][1] <= 20'h7ffff;
            tmp[240][0][1] <= 20'h00000;
            tmp[241][0][1] <= 20'h00000;
            tmp[242][0][1] <= 20'h00000;
            tmp[243][0][1] <= 20'h7ffff;
            tmp[244][0][1] <= 20'h00000;
            tmp[245][0][1] <= 20'h7ffff;
            tmp[246][0][1] <= 20'h7ffff;
            tmp[247][0][1] <= 20'h7ffff;
            tmp[248][0][1] <= 20'h00000;
            tmp[249][0][1] <= 20'h7ffff;
            tmp[250][0][1] <= 20'h7ffff;
            tmp[251][0][1] <= 20'h7ffff;
            tmp[252][0][1] <= 20'h7ffff;
            tmp[253][0][1] <= 20'h7ffff;
            tmp[254][0][1] <= 20'h7ffff;
            tmp[255][0][1] <= 20'h7ffff;
            tmp[256][0][1] <= 20'h00000;
            tmp[257][0][1] <= 20'h00000;
            tmp[258][0][1] <= 20'h00000;
            tmp[259][0][1] <= 20'h00000;
            tmp[260][0][1] <= 20'h00000;
            tmp[261][0][1] <= 20'h00000;
            tmp[262][0][1] <= 20'h00000;
            tmp[263][0][1] <= 20'h7ffff;
            tmp[264][0][1] <= 20'h00000;
            tmp[265][0][1] <= 20'h00000;
            tmp[266][0][1] <= 20'h00000;
            tmp[267][0][1] <= 20'h00000;
            tmp[268][0][1] <= 20'h00000;
            tmp[269][0][1] <= 20'h00000;
            tmp[270][0][1] <= 20'h00000;
            tmp[271][0][1] <= 20'h7ffff;
            tmp[272][0][1] <= 20'h00000;
            tmp[273][0][1] <= 20'h00000;
            tmp[274][0][1] <= 20'h00000;
            tmp[275][0][1] <= 20'h00000;
            tmp[276][0][1] <= 20'h00000;
            tmp[277][0][1] <= 20'h00000;
            tmp[278][0][1] <= 20'h00000;
            tmp[279][0][1] <= 20'h7ffff;
            tmp[280][0][1] <= 20'h00000;
            tmp[281][0][1] <= 20'h00000;
            tmp[282][0][1] <= 20'h00000;
            tmp[283][0][1] <= 20'h7ffff;
            tmp[284][0][1] <= 20'h00000;
            tmp[285][0][1] <= 20'h7ffff;
            tmp[286][0][1] <= 20'h7ffff;
            tmp[287][0][1] <= 20'h7ffff;
            tmp[288][0][1] <= 20'h00000;
            tmp[289][0][1] <= 20'h00000;
            tmp[290][0][1] <= 20'h00000;
            tmp[291][0][1] <= 20'h00000;
            tmp[292][0][1] <= 20'h00000;
            tmp[293][0][1] <= 20'h00000;
            tmp[294][0][1] <= 20'h00000;
            tmp[295][0][1] <= 20'h7ffff;
            tmp[296][0][1] <= 20'h00000;
            tmp[297][0][1] <= 20'h00000;
            tmp[298][0][1] <= 20'h00000;
            tmp[299][0][1] <= 20'h7ffff;
            tmp[300][0][1] <= 20'h00000;
            tmp[301][0][1] <= 20'h7ffff;
            tmp[302][0][1] <= 20'h7ffff;
            tmp[303][0][1] <= 20'h7ffff;
            tmp[304][0][1] <= 20'h00000;
            tmp[305][0][1] <= 20'h00000;
            tmp[306][0][1] <= 20'h00000;
            tmp[307][0][1] <= 20'h7ffff;
            tmp[308][0][1] <= 20'h00000;
            tmp[309][0][1] <= 20'h7ffff;
            tmp[310][0][1] <= 20'h7ffff;
            tmp[311][0][1] <= 20'h7ffff;
            tmp[312][0][1] <= 20'h00000;
            tmp[313][0][1] <= 20'h7ffff;
            tmp[314][0][1] <= 20'h7ffff;
            tmp[315][0][1] <= 20'h7ffff;
            tmp[316][0][1] <= 20'h00000;
            tmp[317][0][1] <= 20'h7ffff;
            tmp[318][0][1] <= 20'h7ffff;
            tmp[319][0][1] <= 20'h7ffff;
            tmp[320][0][1] <= 20'h00000;
            tmp[321][0][1] <= 20'h00000;
            tmp[322][0][1] <= 20'h00000;
            tmp[323][0][1] <= 20'h00000;
            tmp[324][0][1] <= 20'h00000;
            tmp[325][0][1] <= 20'h00000;
            tmp[326][0][1] <= 20'h00000;
            tmp[327][0][1] <= 20'h7ffff;
            tmp[328][0][1] <= 20'h00000;
            tmp[329][0][1] <= 20'h00000;
            tmp[330][0][1] <= 20'h00000;
            tmp[331][0][1] <= 20'h7ffff;
            tmp[332][0][1] <= 20'h00000;
            tmp[333][0][1] <= 20'h7ffff;
            tmp[334][0][1] <= 20'h7ffff;
            tmp[335][0][1] <= 20'h7ffff;
            tmp[336][0][1] <= 20'h00000;
            tmp[337][0][1] <= 20'h00000;
            tmp[338][0][1] <= 20'h00000;
            tmp[339][0][1] <= 20'h7ffff;
            tmp[340][0][1] <= 20'h00000;
            tmp[341][0][1] <= 20'h7ffff;
            tmp[342][0][1] <= 20'h7ffff;
            tmp[343][0][1] <= 20'h7ffff;
            tmp[344][0][1] <= 20'h00000;
            tmp[345][0][1] <= 20'h7ffff;
            tmp[346][0][1] <= 20'h00000;
            tmp[347][0][1] <= 20'h7ffff;
            tmp[348][0][1] <= 20'h00000;
            tmp[349][0][1] <= 20'h7ffff;
            tmp[350][0][1] <= 20'h7ffff;
            tmp[351][0][1] <= 20'h7ffff;
            tmp[352][0][1] <= 20'h00000;
            tmp[353][0][1] <= 20'h00000;
            tmp[354][0][1] <= 20'h00000;
            tmp[355][0][1] <= 20'h7ffff;
            tmp[356][0][1] <= 20'h00000;
            tmp[357][0][1] <= 20'h7ffff;
            tmp[358][0][1] <= 20'h00000;
            tmp[359][0][1] <= 20'h7ffff;
            tmp[360][0][1] <= 20'h00000;
            tmp[361][0][1] <= 20'h7ffff;
            tmp[362][0][1] <= 20'h00000;
            tmp[363][0][1] <= 20'h7ffff;
            tmp[364][0][1] <= 20'h00000;
            tmp[365][0][1] <= 20'h7ffff;
            tmp[366][0][1] <= 20'h7ffff;
            tmp[367][0][1] <= 20'h7ffff;
            tmp[368][0][1] <= 20'h00000;
            tmp[369][0][1] <= 20'h00000;
            tmp[370][0][1] <= 20'h00000;
            tmp[371][0][1] <= 20'h7ffff;
            tmp[372][0][1] <= 20'h00000;
            tmp[373][0][1] <= 20'h7ffff;
            tmp[374][0][1] <= 20'h7ffff;
            tmp[375][0][1] <= 20'h7ffff;
            tmp[376][0][1] <= 20'h00000;
            tmp[377][0][1] <= 20'h7ffff;
            tmp[378][0][1] <= 20'h7ffff;
            tmp[379][0][1] <= 20'h7ffff;
            tmp[380][0][1] <= 20'h7ffff;
            tmp[381][0][1] <= 20'h7ffff;
            tmp[382][0][1] <= 20'h7ffff;
            tmp[383][0][1] <= 20'h7ffff;
            tmp[384][0][1] <= 20'h00000;
            tmp[385][0][1] <= 20'h00000;
            tmp[386][0][1] <= 20'h00000;
            tmp[387][0][1] <= 20'h00000;
            tmp[388][0][1] <= 20'h00000;
            tmp[389][0][1] <= 20'h00000;
            tmp[390][0][1] <= 20'h00000;
            tmp[391][0][1] <= 20'h7ffff;
            tmp[392][0][1] <= 20'h00000;
            tmp[393][0][1] <= 20'h00000;
            tmp[394][0][1] <= 20'h00000;
            tmp[395][0][1] <= 20'h7ffff;
            tmp[396][0][1] <= 20'h00000;
            tmp[397][0][1] <= 20'h7ffff;
            tmp[398][0][1] <= 20'h7ffff;
            tmp[399][0][1] <= 20'h7ffff;
            tmp[400][0][1] <= 20'h00000;
            tmp[401][0][1] <= 20'h00000;
            tmp[402][0][1] <= 20'h00000;
            tmp[403][0][1] <= 20'h7ffff;
            tmp[404][0][1] <= 20'h00000;
            tmp[405][0][1] <= 20'h7ffff;
            tmp[406][0][1] <= 20'h7ffff;
            tmp[407][0][1] <= 20'h7ffff;
            tmp[408][0][1] <= 20'h00000;
            tmp[409][0][1] <= 20'h7ffff;
            tmp[410][0][1] <= 20'h00000;
            tmp[411][0][1] <= 20'h7ffff;
            tmp[412][0][1] <= 20'h00000;
            tmp[413][0][1] <= 20'h7ffff;
            tmp[414][0][1] <= 20'h7ffff;
            tmp[415][0][1] <= 20'h7ffff;
            tmp[416][0][1] <= 20'h00000;
            tmp[417][0][1] <= 20'h00000;
            tmp[418][0][1] <= 20'h00000;
            tmp[419][0][1] <= 20'h7ffff;
            tmp[420][0][1] <= 20'h00000;
            tmp[421][0][1] <= 20'h7ffff;
            tmp[422][0][1] <= 20'h00000;
            tmp[423][0][1] <= 20'h7ffff;
            tmp[424][0][1] <= 20'h00000;
            tmp[425][0][1] <= 20'h7ffff;
            tmp[426][0][1] <= 20'h00000;
            tmp[427][0][1] <= 20'h7ffff;
            tmp[428][0][1] <= 20'h00000;
            tmp[429][0][1] <= 20'h7ffff;
            tmp[430][0][1] <= 20'h7ffff;
            tmp[431][0][1] <= 20'h7ffff;
            tmp[432][0][1] <= 20'h00000;
            tmp[433][0][1] <= 20'h00000;
            tmp[434][0][1] <= 20'h00000;
            tmp[435][0][1] <= 20'h7ffff;
            tmp[436][0][1] <= 20'h00000;
            tmp[437][0][1] <= 20'h7ffff;
            tmp[438][0][1] <= 20'h7ffff;
            tmp[439][0][1] <= 20'h7ffff;
            tmp[440][0][1] <= 20'h00000;
            tmp[441][0][1] <= 20'h7ffff;
            tmp[442][0][1] <= 20'h7ffff;
            tmp[443][0][1] <= 20'h7ffff;
            tmp[444][0][1] <= 20'h7ffff;
            tmp[445][0][1] <= 20'h7ffff;
            tmp[446][0][1] <= 20'h7ffff;
            tmp[447][0][1] <= 20'h7ffff;
            tmp[448][0][1] <= 20'h00000;
            tmp[449][0][1] <= 20'h00000;
            tmp[450][0][1] <= 20'h00000;
            tmp[451][0][1] <= 20'h7ffff;
            tmp[452][0][1] <= 20'h00000;
            tmp[453][0][1] <= 20'h7ffff;
            tmp[454][0][1] <= 20'h00000;
            tmp[455][0][1] <= 20'h7ffff;
            tmp[456][0][1] <= 20'h00000;
            tmp[457][0][1] <= 20'h00000;
            tmp[458][0][1] <= 20'h00000;
            tmp[459][0][1] <= 20'h7ffff;
            tmp[460][0][1] <= 20'h00000;
            tmp[461][0][1] <= 20'h7ffff;
            tmp[462][0][1] <= 20'h7ffff;
            tmp[463][0][1] <= 20'h7ffff;
            tmp[464][0][1] <= 20'h00000;
            tmp[465][0][1] <= 20'h00000;
            tmp[466][0][1] <= 20'h00000;
            tmp[467][0][1] <= 20'h7ffff;
            tmp[468][0][1] <= 20'h00000;
            tmp[469][0][1] <= 20'h7ffff;
            tmp[470][0][1] <= 20'h7ffff;
            tmp[471][0][1] <= 20'h7ffff;
            tmp[472][0][1] <= 20'h00000;
            tmp[473][0][1] <= 20'h7ffff;
            tmp[474][0][1] <= 20'h7ffff;
            tmp[475][0][1] <= 20'h7ffff;
            tmp[476][0][1] <= 20'h7ffff;
            tmp[477][0][1] <= 20'h7ffff;
            tmp[478][0][1] <= 20'h7ffff;
            tmp[479][0][1] <= 20'h7ffff;
            tmp[480][0][1] <= 20'h00000;
            tmp[481][0][1] <= 20'h00000;
            tmp[482][0][1] <= 20'h00000;
            tmp[483][0][1] <= 20'h7ffff;
            tmp[484][0][1] <= 20'h00000;
            tmp[485][0][1] <= 20'h7ffff;
            tmp[486][0][1] <= 20'h7ffff;
            tmp[487][0][1] <= 20'h7ffff;
            tmp[488][0][1] <= 20'h00000;
            tmp[489][0][1] <= 20'h7ffff;
            tmp[490][0][1] <= 20'h7ffff;
            tmp[491][0][1] <= 20'h7ffff;
            tmp[492][0][1] <= 20'h7ffff;
            tmp[493][0][1] <= 20'h7ffff;
            tmp[494][0][1] <= 20'h7ffff;
            tmp[495][0][1] <= 20'h7ffff;
            tmp[496][0][1] <= 20'h00000;
            tmp[497][0][1] <= 20'h7ffff;
            tmp[498][0][1] <= 20'h7ffff;
            tmp[499][0][1] <= 20'h7ffff;
            tmp[500][0][1] <= 20'h00000;
            tmp[501][0][1] <= 20'h7ffff;
            tmp[502][0][1] <= 20'h7ffff;
            tmp[503][0][1] <= 20'h7ffff;
            tmp[504][0][1] <= 20'h00000;
            tmp[505][0][1] <= 20'h7ffff;
            tmp[506][0][1] <= 20'h7ffff;
            tmp[507][0][1] <= 20'h7ffff;
            tmp[508][0][1] <= 20'h7ffff;
            tmp[509][0][1] <= 20'h7ffff;
            tmp[510][0][1] <= 20'h7ffff;
            tmp[511][0][1] <= 20'h7ffff;
            tmp[512][0][1] <= 20'h00000;
            tmp[513][0][1] <= 20'h00000;
            tmp[514][0][1] <= 20'h00000;
            tmp[515][0][1] <= 20'h00000;
            tmp[516][0][1] <= 20'h00000;
            tmp[517][0][1] <= 20'h00000;
            tmp[518][0][1] <= 20'h00000;
            tmp[519][0][1] <= 20'h7ffff;
            tmp[520][0][1] <= 20'h00000;
            tmp[521][0][1] <= 20'h00000;
            tmp[522][0][1] <= 20'h00000;
            tmp[523][0][1] <= 20'h00000;
            tmp[524][0][1] <= 20'h00000;
            tmp[525][0][1] <= 20'h00000;
            tmp[526][0][1] <= 20'h00000;
            tmp[527][0][1] <= 20'h7ffff;
            tmp[528][0][1] <= 20'h00000;
            tmp[529][0][1] <= 20'h00000;
            tmp[530][0][1] <= 20'h00000;
            tmp[531][0][1] <= 20'h00000;
            tmp[532][0][1] <= 20'h00000;
            tmp[533][0][1] <= 20'h00000;
            tmp[534][0][1] <= 20'h00000;
            tmp[535][0][1] <= 20'h7ffff;
            tmp[536][0][1] <= 20'h00000;
            tmp[537][0][1] <= 20'h00000;
            tmp[538][0][1] <= 20'h00000;
            tmp[539][0][1] <= 20'h7ffff;
            tmp[540][0][1] <= 20'h00000;
            tmp[541][0][1] <= 20'h7ffff;
            tmp[542][0][1] <= 20'h7ffff;
            tmp[543][0][1] <= 20'h7ffff;
            tmp[544][0][1] <= 20'h00000;
            tmp[545][0][1] <= 20'h00000;
            tmp[546][0][1] <= 20'h00000;
            tmp[547][0][1] <= 20'h00000;
            tmp[548][0][1] <= 20'h00000;
            tmp[549][0][1] <= 20'h00000;
            tmp[550][0][1] <= 20'h00000;
            tmp[551][0][1] <= 20'h7ffff;
            tmp[552][0][1] <= 20'h00000;
            tmp[553][0][1] <= 20'h00000;
            tmp[554][0][1] <= 20'h00000;
            tmp[555][0][1] <= 20'h7ffff;
            tmp[556][0][1] <= 20'h00000;
            tmp[557][0][1] <= 20'h7ffff;
            tmp[558][0][1] <= 20'h7ffff;
            tmp[559][0][1] <= 20'h7ffff;
            tmp[560][0][1] <= 20'h00000;
            tmp[561][0][1] <= 20'h00000;
            tmp[562][0][1] <= 20'h00000;
            tmp[563][0][1] <= 20'h7ffff;
            tmp[564][0][1] <= 20'h00000;
            tmp[565][0][1] <= 20'h7ffff;
            tmp[566][0][1] <= 20'h7ffff;
            tmp[567][0][1] <= 20'h7ffff;
            tmp[568][0][1] <= 20'h00000;
            tmp[569][0][1] <= 20'h7ffff;
            tmp[570][0][1] <= 20'h00000;
            tmp[571][0][1] <= 20'h7ffff;
            tmp[572][0][1] <= 20'h00000;
            tmp[573][0][1] <= 20'h7ffff;
            tmp[574][0][1] <= 20'h7ffff;
            tmp[575][0][1] <= 20'h7ffff;
            tmp[576][0][1] <= 20'h00000;
            tmp[577][0][1] <= 20'h00000;
            tmp[578][0][1] <= 20'h00000;
            tmp[579][0][1] <= 20'h00000;
            tmp[580][0][1] <= 20'h00000;
            tmp[581][0][1] <= 20'h00000;
            tmp[582][0][1] <= 20'h00000;
            tmp[583][0][1] <= 20'h7ffff;
            tmp[584][0][1] <= 20'h00000;
            tmp[585][0][1] <= 20'h00000;
            tmp[586][0][1] <= 20'h00000;
            tmp[587][0][1] <= 20'h7ffff;
            tmp[588][0][1] <= 20'h00000;
            tmp[589][0][1] <= 20'h7ffff;
            tmp[590][0][1] <= 20'h7ffff;
            tmp[591][0][1] <= 20'h7ffff;
            tmp[592][0][1] <= 20'h00000;
            tmp[593][0][1] <= 20'h00000;
            tmp[594][0][1] <= 20'h00000;
            tmp[595][0][1] <= 20'h7ffff;
            tmp[596][0][1] <= 20'h00000;
            tmp[597][0][1] <= 20'h7ffff;
            tmp[598][0][1] <= 20'h7ffff;
            tmp[599][0][1] <= 20'h7ffff;
            tmp[600][0][1] <= 20'h00000;
            tmp[601][0][1] <= 20'h7ffff;
            tmp[602][0][1] <= 20'h00000;
            tmp[603][0][1] <= 20'h7ffff;
            tmp[604][0][1] <= 20'h00000;
            tmp[605][0][1] <= 20'h7ffff;
            tmp[606][0][1] <= 20'h7ffff;
            tmp[607][0][1] <= 20'h7ffff;
            tmp[608][0][1] <= 20'h00000;
            tmp[609][0][1] <= 20'h00000;
            tmp[610][0][1] <= 20'h00000;
            tmp[611][0][1] <= 20'h7ffff;
            tmp[612][0][1] <= 20'h00000;
            tmp[613][0][1] <= 20'h7ffff;
            tmp[614][0][1] <= 20'h00000;
            tmp[615][0][1] <= 20'h7ffff;
            tmp[616][0][1] <= 20'h00000;
            tmp[617][0][1] <= 20'h7ffff;
            tmp[618][0][1] <= 20'h00000;
            tmp[619][0][1] <= 20'h7ffff;
            tmp[620][0][1] <= 20'h00000;
            tmp[621][0][1] <= 20'h7ffff;
            tmp[622][0][1] <= 20'h7ffff;
            tmp[623][0][1] <= 20'h7ffff;
            tmp[624][0][1] <= 20'h00000;
            tmp[625][0][1] <= 20'h00000;
            tmp[626][0][1] <= 20'h00000;
            tmp[627][0][1] <= 20'h7ffff;
            tmp[628][0][1] <= 20'h00000;
            tmp[629][0][1] <= 20'h7ffff;
            tmp[630][0][1] <= 20'h7ffff;
            tmp[631][0][1] <= 20'h7ffff;
            tmp[632][0][1] <= 20'h00000;
            tmp[633][0][1] <= 20'h7ffff;
            tmp[634][0][1] <= 20'h7ffff;
            tmp[635][0][1] <= 20'h7ffff;
            tmp[636][0][1] <= 20'h7ffff;
            tmp[637][0][1] <= 20'h7ffff;
            tmp[638][0][1] <= 20'h7ffff;
            tmp[639][0][1] <= 20'h7ffff;
            tmp[640][0][1] <= 20'h00000;
            tmp[641][0][1] <= 20'h00000;
            tmp[642][0][1] <= 20'h00000;
            tmp[643][0][1] <= 20'h00000;
            tmp[644][0][1] <= 20'h00000;
            tmp[645][0][1] <= 20'h00000;
            tmp[646][0][1] <= 20'h00000;
            tmp[647][0][1] <= 20'h7ffff;
            tmp[648][0][1] <= 20'h00000;
            tmp[649][0][1] <= 20'h00000;
            tmp[650][0][1] <= 20'h00000;
            tmp[651][0][1] <= 20'h7ffff;
            tmp[652][0][1] <= 20'h00000;
            tmp[653][0][1] <= 20'h7ffff;
            tmp[654][0][1] <= 20'h7ffff;
            tmp[655][0][1] <= 20'h7ffff;
            tmp[656][0][1] <= 20'h00000;
            tmp[657][0][1] <= 20'h00000;
            tmp[658][0][1] <= 20'h00000;
            tmp[659][0][1] <= 20'h7ffff;
            tmp[660][0][1] <= 20'h00000;
            tmp[661][0][1] <= 20'h7ffff;
            tmp[662][0][1] <= 20'h7ffff;
            tmp[663][0][1] <= 20'h7ffff;
            tmp[664][0][1] <= 20'h00000;
            tmp[665][0][1] <= 20'h7ffff;
            tmp[666][0][1] <= 20'h00000;
            tmp[667][0][1] <= 20'h7ffff;
            tmp[668][0][1] <= 20'h00000;
            tmp[669][0][1] <= 20'h7ffff;
            tmp[670][0][1] <= 20'h7ffff;
            tmp[671][0][1] <= 20'h7ffff;
            tmp[672][0][1] <= 20'h00000;
            tmp[673][0][1] <= 20'h00000;
            tmp[674][0][1] <= 20'h00000;
            tmp[675][0][1] <= 20'h7ffff;
            tmp[676][0][1] <= 20'h00000;
            tmp[677][0][1] <= 20'h7ffff;
            tmp[678][0][1] <= 20'h00000;
            tmp[679][0][1] <= 20'h7ffff;
            tmp[680][0][1] <= 20'h00000;
            tmp[681][0][1] <= 20'h00000;
            tmp[682][0][1] <= 20'h00000;
            tmp[683][0][1] <= 20'h7ffff;
            tmp[684][0][1] <= 20'h00000;
            tmp[685][0][1] <= 20'h7ffff;
            tmp[686][0][1] <= 20'h7ffff;
            tmp[687][0][1] <= 20'h7ffff;
            tmp[688][0][1] <= 20'h00000;
            tmp[689][0][1] <= 20'h00000;
            tmp[690][0][1] <= 20'h00000;
            tmp[691][0][1] <= 20'h7ffff;
            tmp[692][0][1] <= 20'h00000;
            tmp[693][0][1] <= 20'h7ffff;
            tmp[694][0][1] <= 20'h7ffff;
            tmp[695][0][1] <= 20'h7ffff;
            tmp[696][0][1] <= 20'h00000;
            tmp[697][0][1] <= 20'h7ffff;
            tmp[698][0][1] <= 20'h7ffff;
            tmp[699][0][1] <= 20'h7ffff;
            tmp[700][0][1] <= 20'h7ffff;
            tmp[701][0][1] <= 20'h7ffff;
            tmp[702][0][1] <= 20'h7ffff;
            tmp[703][0][1] <= 20'h7ffff;
            tmp[704][0][1] <= 20'h00000;
            tmp[705][0][1] <= 20'h00000;
            tmp[706][0][1] <= 20'h00000;
            tmp[707][0][1] <= 20'h7ffff;
            tmp[708][0][1] <= 20'h00000;
            tmp[709][0][1] <= 20'h7ffff;
            tmp[710][0][1] <= 20'h00000;
            tmp[711][0][1] <= 20'h7ffff;
            tmp[712][0][1] <= 20'h00000;
            tmp[713][0][1] <= 20'h00000;
            tmp[714][0][1] <= 20'h00000;
            tmp[715][0][1] <= 20'h7ffff;
            tmp[716][0][1] <= 20'h00000;
            tmp[717][0][1] <= 20'h7ffff;
            tmp[718][0][1] <= 20'h7ffff;
            tmp[719][0][1] <= 20'h7ffff;
            tmp[720][0][1] <= 20'h00000;
            tmp[721][0][1] <= 20'h00000;
            tmp[722][0][1] <= 20'h00000;
            tmp[723][0][1] <= 20'h7ffff;
            tmp[724][0][1] <= 20'h00000;
            tmp[725][0][1] <= 20'h7ffff;
            tmp[726][0][1] <= 20'h7ffff;
            tmp[727][0][1] <= 20'h7ffff;
            tmp[728][0][1] <= 20'h00000;
            tmp[729][0][1] <= 20'h7ffff;
            tmp[730][0][1] <= 20'h7ffff;
            tmp[731][0][1] <= 20'h7ffff;
            tmp[732][0][1] <= 20'h7ffff;
            tmp[733][0][1] <= 20'h7ffff;
            tmp[734][0][1] <= 20'h7ffff;
            tmp[735][0][1] <= 20'h7ffff;
            tmp[736][0][1] <= 20'h00000;
            tmp[737][0][1] <= 20'h00000;
            tmp[738][0][1] <= 20'h00000;
            tmp[739][0][1] <= 20'h7ffff;
            tmp[740][0][1] <= 20'h00000;
            tmp[741][0][1] <= 20'h7ffff;
            tmp[742][0][1] <= 20'h7ffff;
            tmp[743][0][1] <= 20'h7ffff;
            tmp[744][0][1] <= 20'h00000;
            tmp[745][0][1] <= 20'h7ffff;
            tmp[746][0][1] <= 20'h7ffff;
            tmp[747][0][1] <= 20'h7ffff;
            tmp[748][0][1] <= 20'h7ffff;
            tmp[749][0][1] <= 20'h7ffff;
            tmp[750][0][1] <= 20'h7ffff;
            tmp[751][0][1] <= 20'h7ffff;
            tmp[752][0][1] <= 20'h00000;
            tmp[753][0][1] <= 20'h7ffff;
            tmp[754][0][1] <= 20'h7ffff;
            tmp[755][0][1] <= 20'h7ffff;
            tmp[756][0][1] <= 20'h00000;
            tmp[757][0][1] <= 20'h7ffff;
            tmp[758][0][1] <= 20'h7ffff;
            tmp[759][0][1] <= 20'h7ffff;
            tmp[760][0][1] <= 20'h00000;
            tmp[761][0][1] <= 20'h7ffff;
            tmp[762][0][1] <= 20'h7ffff;
            tmp[763][0][1] <= 20'h7ffff;
            tmp[764][0][1] <= 20'h7ffff;
            tmp[765][0][1] <= 20'h7ffff;
            tmp[766][0][1] <= 20'h7ffff;
            tmp[767][0][1] <= 20'h7ffff;
            tmp[768][0][1] <= 20'h00000;
            tmp[769][0][1] <= 20'h00000;
            tmp[770][0][1] <= 20'h00000;
            tmp[771][0][1] <= 20'h00000;
            tmp[772][0][1] <= 20'h00000;
            tmp[773][0][1] <= 20'h00000;
            tmp[774][0][1] <= 20'h00000;
            tmp[775][0][1] <= 20'h7ffff;
            tmp[776][0][1] <= 20'h00000;
            tmp[777][0][1] <= 20'h00000;
            tmp[778][0][1] <= 20'h00000;
            tmp[779][0][1] <= 20'h7ffff;
            tmp[780][0][1] <= 20'h00000;
            tmp[781][0][1] <= 20'h7ffff;
            tmp[782][0][1] <= 20'h7ffff;
            tmp[783][0][1] <= 20'h7ffff;
            tmp[784][0][1] <= 20'h00000;
            tmp[785][0][1] <= 20'h00000;
            tmp[786][0][1] <= 20'h00000;
            tmp[787][0][1] <= 20'h7ffff;
            tmp[788][0][1] <= 20'h00000;
            tmp[789][0][1] <= 20'h7ffff;
            tmp[790][0][1] <= 20'h00000;
            tmp[791][0][1] <= 20'h7ffff;
            tmp[792][0][1] <= 20'h00000;
            tmp[793][0][1] <= 20'h7ffff;
            tmp[794][0][1] <= 20'h00000;
            tmp[795][0][1] <= 20'h7ffff;
            tmp[796][0][1] <= 20'h00000;
            tmp[797][0][1] <= 20'h7ffff;
            tmp[798][0][1] <= 20'h7ffff;
            tmp[799][0][1] <= 20'h7ffff;
            tmp[800][0][1] <= 20'h00000;
            tmp[801][0][1] <= 20'h00000;
            tmp[802][0][1] <= 20'h00000;
            tmp[803][0][1] <= 20'h7ffff;
            tmp[804][0][1] <= 20'h00000;
            tmp[805][0][1] <= 20'h7ffff;
            tmp[806][0][1] <= 20'h00000;
            tmp[807][0][1] <= 20'h7ffff;
            tmp[808][0][1] <= 20'h00000;
            tmp[809][0][1] <= 20'h00000;
            tmp[810][0][1] <= 20'h00000;
            tmp[811][0][1] <= 20'h7ffff;
            tmp[812][0][1] <= 20'h00000;
            tmp[813][0][1] <= 20'h7ffff;
            tmp[814][0][1] <= 20'h7ffff;
            tmp[815][0][1] <= 20'h7ffff;
            tmp[816][0][1] <= 20'h00000;
            tmp[817][0][1] <= 20'h00000;
            tmp[818][0][1] <= 20'h00000;
            tmp[819][0][1] <= 20'h7ffff;
            tmp[820][0][1] <= 20'h00000;
            tmp[821][0][1] <= 20'h7ffff;
            tmp[822][0][1] <= 20'h7ffff;
            tmp[823][0][1] <= 20'h7ffff;
            tmp[824][0][1] <= 20'h00000;
            tmp[825][0][1] <= 20'h7ffff;
            tmp[826][0][1] <= 20'h7ffff;
            tmp[827][0][1] <= 20'h7ffff;
            tmp[828][0][1] <= 20'h7ffff;
            tmp[829][0][1] <= 20'h7ffff;
            tmp[830][0][1] <= 20'h7ffff;
            tmp[831][0][1] <= 20'h7ffff;
            tmp[832][0][1] <= 20'h00000;
            tmp[833][0][1] <= 20'h00000;
            tmp[834][0][1] <= 20'h00000;
            tmp[835][0][1] <= 20'h7ffff;
            tmp[836][0][1] <= 20'h00000;
            tmp[837][0][1] <= 20'h00000;
            tmp[838][0][1] <= 20'h00000;
            tmp[839][0][1] <= 20'h7ffff;
            tmp[840][0][1] <= 20'h00000;
            tmp[841][0][1] <= 20'h00000;
            tmp[842][0][1] <= 20'h00000;
            tmp[843][0][1] <= 20'h7ffff;
            tmp[844][0][1] <= 20'h00000;
            tmp[845][0][1] <= 20'h7ffff;
            tmp[846][0][1] <= 20'h7ffff;
            tmp[847][0][1] <= 20'h7ffff;
            tmp[848][0][1] <= 20'h00000;
            tmp[849][0][1] <= 20'h00000;
            tmp[850][0][1] <= 20'h00000;
            tmp[851][0][1] <= 20'h7ffff;
            tmp[852][0][1] <= 20'h00000;
            tmp[853][0][1] <= 20'h7ffff;
            tmp[854][0][1] <= 20'h7ffff;
            tmp[855][0][1] <= 20'h7ffff;
            tmp[856][0][1] <= 20'h00000;
            tmp[857][0][1] <= 20'h7ffff;
            tmp[858][0][1] <= 20'h7ffff;
            tmp[859][0][1] <= 20'h7ffff;
            tmp[860][0][1] <= 20'h7ffff;
            tmp[861][0][1] <= 20'h7ffff;
            tmp[862][0][1] <= 20'h7ffff;
            tmp[863][0][1] <= 20'h7ffff;
            tmp[864][0][1] <= 20'h00000;
            tmp[865][0][1] <= 20'h00000;
            tmp[866][0][1] <= 20'h00000;
            tmp[867][0][1] <= 20'h7ffff;
            tmp[868][0][1] <= 20'h00000;
            tmp[869][0][1] <= 20'h7ffff;
            tmp[870][0][1] <= 20'h7ffff;
            tmp[871][0][1] <= 20'h7ffff;
            tmp[872][0][1] <= 20'h00000;
            tmp[873][0][1] <= 20'h7ffff;
            tmp[874][0][1] <= 20'h7ffff;
            tmp[875][0][1] <= 20'h7ffff;
            tmp[876][0][1] <= 20'h7ffff;
            tmp[877][0][1] <= 20'h7ffff;
            tmp[878][0][1] <= 20'h7ffff;
            tmp[879][0][1] <= 20'h7ffff;
            tmp[880][0][1] <= 20'h00000;
            tmp[881][0][1] <= 20'h7ffff;
            tmp[882][0][1] <= 20'h7ffff;
            tmp[883][0][1] <= 20'h7ffff;
            tmp[884][0][1] <= 20'h00000;
            tmp[885][0][1] <= 20'h7ffff;
            tmp[886][0][1] <= 20'h7ffff;
            tmp[887][0][1] <= 20'h7ffff;
            tmp[888][0][1] <= 20'h00000;
            tmp[889][0][1] <= 20'h7ffff;
            tmp[890][0][1] <= 20'h7ffff;
            tmp[891][0][1] <= 20'h7ffff;
            tmp[892][0][1] <= 20'h7ffff;
            tmp[893][0][1] <= 20'h7ffff;
            tmp[894][0][1] <= 20'h7ffff;
            tmp[895][0][1] <= 20'h7ffff;
            tmp[896][0][1] <= 20'h00000;
            tmp[897][0][1] <= 20'h00000;
            tmp[898][0][1] <= 20'h00000;
            tmp[899][0][1] <= 20'h7ffff;
            tmp[900][0][1] <= 20'h00000;
            tmp[901][0][1] <= 20'h00000;
            tmp[902][0][1] <= 20'h00000;
            tmp[903][0][1] <= 20'h7ffff;
            tmp[904][0][1] <= 20'h00000;
            tmp[905][0][1] <= 20'h00000;
            tmp[906][0][1] <= 20'h00000;
            tmp[907][0][1] <= 20'h7ffff;
            tmp[908][0][1] <= 20'h00000;
            tmp[909][0][1] <= 20'h7ffff;
            tmp[910][0][1] <= 20'h7ffff;
            tmp[911][0][1] <= 20'h7ffff;
            tmp[912][0][1] <= 20'h00000;
            tmp[913][0][1] <= 20'h00000;
            tmp[914][0][1] <= 20'h00000;
            tmp[915][0][1] <= 20'h7ffff;
            tmp[916][0][1] <= 20'h00000;
            tmp[917][0][1] <= 20'h7ffff;
            tmp[918][0][1] <= 20'h7ffff;
            tmp[919][0][1] <= 20'h7ffff;
            tmp[920][0][1] <= 20'h00000;
            tmp[921][0][1] <= 20'h7ffff;
            tmp[922][0][1] <= 20'h7ffff;
            tmp[923][0][1] <= 20'h7ffff;
            tmp[924][0][1] <= 20'h7ffff;
            tmp[925][0][1] <= 20'h7ffff;
            tmp[926][0][1] <= 20'h7ffff;
            tmp[927][0][1] <= 20'h7ffff;
            tmp[928][0][1] <= 20'h00000;
            tmp[929][0][1] <= 20'h00000;
            tmp[930][0][1] <= 20'h00000;
            tmp[931][0][1] <= 20'h7ffff;
            tmp[932][0][1] <= 20'h00000;
            tmp[933][0][1] <= 20'h7ffff;
            tmp[934][0][1] <= 20'h7ffff;
            tmp[935][0][1] <= 20'h7ffff;
            tmp[936][0][1] <= 20'h00000;
            tmp[937][0][1] <= 20'h7ffff;
            tmp[938][0][1] <= 20'h7ffff;
            tmp[939][0][1] <= 20'h7ffff;
            tmp[940][0][1] <= 20'h00000;
            tmp[941][0][1] <= 20'h7ffff;
            tmp[942][0][1] <= 20'h7ffff;
            tmp[943][0][1] <= 20'h7ffff;
            tmp[944][0][1] <= 20'h00000;
            tmp[945][0][1] <= 20'h7ffff;
            tmp[946][0][1] <= 20'h7ffff;
            tmp[947][0][1] <= 20'h7ffff;
            tmp[948][0][1] <= 20'h00000;
            tmp[949][0][1] <= 20'h7ffff;
            tmp[950][0][1] <= 20'h7ffff;
            tmp[951][0][1] <= 20'h7ffff;
            tmp[952][0][1] <= 20'h00000;
            tmp[953][0][1] <= 20'h7ffff;
            tmp[954][0][1] <= 20'h7ffff;
            tmp[955][0][1] <= 20'h7ffff;
            tmp[956][0][1] <= 20'h7ffff;
            tmp[957][0][1] <= 20'h7ffff;
            tmp[958][0][1] <= 20'h7ffff;
            tmp[959][0][1] <= 20'h7ffff;
            tmp[960][0][1] <= 20'h00000;
            tmp[961][0][1] <= 20'h00000;
            tmp[962][0][1] <= 20'h00000;
            tmp[963][0][1] <= 20'h7ffff;
            tmp[964][0][1] <= 20'h00000;
            tmp[965][0][1] <= 20'h7ffff;
            tmp[966][0][1] <= 20'h7ffff;
            tmp[967][0][1] <= 20'h7ffff;
            tmp[968][0][1] <= 20'h00000;
            tmp[969][0][1] <= 20'h7ffff;
            tmp[970][0][1] <= 20'h7ffff;
            tmp[971][0][1] <= 20'h7ffff;
            tmp[972][0][1] <= 20'h00000;
            tmp[973][0][1] <= 20'h7ffff;
            tmp[974][0][1] <= 20'h7ffff;
            tmp[975][0][1] <= 20'h7ffff;
            tmp[976][0][1] <= 20'h00000;
            tmp[977][0][1] <= 20'h7ffff;
            tmp[978][0][1] <= 20'h00000;
            tmp[979][0][1] <= 20'h7ffff;
            tmp[980][0][1] <= 20'h00000;
            tmp[981][0][1] <= 20'h7ffff;
            tmp[982][0][1] <= 20'h7ffff;
            tmp[983][0][1] <= 20'h7ffff;
            tmp[984][0][1] <= 20'h00000;
            tmp[985][0][1] <= 20'h7ffff;
            tmp[986][0][1] <= 20'h7ffff;
            tmp[987][0][1] <= 20'h7ffff;
            tmp[988][0][1] <= 20'h7ffff;
            tmp[989][0][1] <= 20'h7ffff;
            tmp[990][0][1] <= 20'h7ffff;
            tmp[991][0][1] <= 20'h7ffff;
            tmp[992][0][1] <= 20'h00000;
            tmp[993][0][1] <= 20'h7ffff;
            tmp[994][0][1] <= 20'h00000;
            tmp[995][0][1] <= 20'h7ffff;
            tmp[996][0][1] <= 20'h00000;
            tmp[997][0][1] <= 20'h7ffff;
            tmp[998][0][1] <= 20'h7ffff;
            tmp[999][0][1] <= 20'h7ffff;
            tmp[1000][0][1] <= 20'h00000;
            tmp[1001][0][1] <= 20'h7ffff;
            tmp[1002][0][1] <= 20'h7ffff;
            tmp[1003][0][1] <= 20'h7ffff;
            tmp[1004][0][1] <= 20'h7ffff;
            tmp[1005][0][1] <= 20'h7ffff;
            tmp[1006][0][1] <= 20'h7ffff;
            tmp[1007][0][1] <= 20'h7ffff;
            tmp[1008][0][1] <= 20'h00000;
            tmp[1009][0][1] <= 20'h7ffff;
            tmp[1010][0][1] <= 20'h7ffff;
            tmp[1011][0][1] <= 20'h7ffff;
            tmp[1012][0][1] <= 20'h7ffff;
            tmp[1013][0][1] <= 20'h7ffff;
            tmp[1014][0][1] <= 20'h7ffff;
            tmp[1015][0][1] <= 20'h7ffff;
            tmp[1016][0][1] <= 20'h7ffff;
            tmp[1017][0][1] <= 20'h7ffff;
            tmp[1018][0][1] <= 20'h7ffff;
            tmp[1019][0][1] <= 20'h7ffff;
            tmp[1020][0][1] <= 20'h7ffff;
            tmp[1021][0][1] <= 20'h7ffff;
            tmp[1022][0][1] <= 20'h7ffff;
            tmp[1023][0][1] <= 20'h7ffff;
        end else begin
            case(stage)
            `DECODE:begin
                done <= 0;
                counter <= counter + 1;
                if (counter >= N-1)begin
                    counter <= 0;
                    stage <= `DONE;
                end else 
                    stage <= stage;

                for (y = 0; y < STEP; y = y + 1)
                    for (x = 0; x < N; x = x + 1)begin
                        tmp[x][y+1][0] <= w[x][y][0];
                    end
            end
            `ENCODE:begin
                done <= 0;
                counter <= counter + 1;
                if(counter >= N-1)begin
                    counter <= 0;
                    stage <= `DECODE;
                    //stage<=`DONE;
                end else 
                    stage <= stage;

                for (y = 0; y < STEP; y = y + 1)
                    for (x = 0; x < N; x = x + 1)begin
                        tmp[x][y+1][1] <= w[x][y][1];
                    end
            end
            default:begin
                done <= 1;
                if(en) 
                    stage <= `ENCODE;
                else 
                    stage <= stage;
            end
            endcase
        end      
    end
endmodule
